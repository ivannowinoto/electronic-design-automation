module sub_module1(
    input wire [2:0] in1,
    input wire [2:0] in2,
    input wire [2:0] in3,
    input wire [2:0] in4,
    input wire [2:0] in5,
    input wire [2:0] in6,
    input wire [2:0] in7,
    input wire [3:0] in8,
    input wire [3:0] in9,
    input wire [3:0] in10,
    input wire [3:0] in11,
    input wire [3:0] in12,
    input wire [3:0] in13,
    input wire [3:0] in14,
    output wire [1:0] out1,
    output wire [1:0] out2,
    output wire [1:0] out3,
    output wire [1:0] out4,
    output wire [1:0] out5,
    output wire [2:0] out6,
    output wire [2:0] out7,
    output wire [2:0] out8,
    output wire [2:0] out9,
    output wire [2:0] out10,
    output wire [3:0] out11,
    output wire [3:0] out12
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
and (w_0208_, w_0701_, w_0639_);
or (w_0648_, w_0332_, w_0578_);
and (w_0219_, in13[2], w_0537_);
and (w_0537_, w_0443_, w_0718_);
or (w_0055_, w_0033_, w_0230_);
not (w_0351_, w_0859_);
not (w_0325_, w_0682_);
and (w_0187_, in1[1], in2[1]);
and (out8[1], w_0394_, w_0174_);
or (out11[3], w_0062_, w_0328_);
and (w_0700_, w_0290_, w_0544_);
or (w_0471_, w_0076_, w_0634_);
or (w_0226_, w_0388_, w_0860_);
and (w_0521_, w_0346_, w_0725_);
or (w_0004_, w_0539_, w_0276_);
not (w_0441_, w_0296_);
or (w_0510_, w_0137_, w_0675_);
not (w_0066_, w_0508_);
or (w_0046_, w_0849_, w_0440_);
and (w_0139_, in3[1], w_0674_);
or (w_0494_, w_0782_, w_0054_);
or (w_0624_, w_0792_, w_0543_);
or (w_0655_, w_0394_, w_0174_);
or (w_0564_, w_0366_, w_0683_);
not (w_0399_, w_0788_);
not (w_0695_, w_0571_);
or (w_0264_, w_0065_, w_0852_);
and (w_0114_, w_0234_, w_0596_);
not (w_0216_, w_0014_);
and (w_0694_, w_0524_, w_0438_);
and (w_0217_, w_0478_, w_0185_);
and (w_0284_, w_0148_, w_0831_);
or (w_0633_, w_0152_, w_0312_);
or (w_0568_, w_0136_, w_0642_);
not (w_0818_, w_0002_);
not (w_0436_, w_0423_);
and (w_0213_, w_0303_, w_0431_);
or (w_0110_, w_0825_, w_0684_);
or (w_0443_, w_0303_, w_0431_);
and (w_0812_, w_0261_, w_0371_);
and (w_0400_, w_0705_, w_0035_);
not (w_0011_, w_0425_);
and (w_0009_, w_0343_, w_0159_);
or (w_0075_, w_0426_, w_0689_);
or (w_0639_, w_0333_, w_0841_);
and (w_0464_, in1[2], w_0336_);
and (w_0278_, in14[3], in8[1]);
or (w_0758_, w_0791_, w_0593_);
or (w_0725_, w_0466_, w_0566_);
or (w_0018_, w_0710_, w_0528_);
and (w_0608_, w_0137_, w_0675_);
or (w_0703_, in13[3], w_0521_);
not (w_0344_, w_0118_);
or (w_0067_, w_0273_, w_0135_);
not (w_0802_, w_0381_);
and (w_0063_, w_0164_, w_0122_);
or (w_0283_, in13[2], w_0537_);
or (w_0589_, in7[1], in2[1]);
or (w_0809_, w_0613_, w_0149_);
and (w_0008_, w_0705_, w_0193_);
and (w_0489_, w_0339_, w_0715_);
and (w_0452_, w_0828_, w_0226_);
or (w_0833_, w_0000_, w_0405_);
and (w_0588_, w_0651_, w_0449_);
or (w_0519_, w_0753_, w_0475_);
or (w_0343_, w_0297_, w_0323_);
or (w_0412_, w_0811_, w_0737_);
and (w_0367_, w_0641_, w_0857_);
and (out12[1], w_0819_, w_0742_);
or (w_0547_, out8[1], w_0401_);
or (w_0415_, w_0729_, w_0848_);
not (w_0222_, in7[2]);
and (w_0375_, in14[2], w_0285_);
or (w_0607_, w_0636_, w_0167_);
and (w_0706_, w_0692_, w_0626_);
and (w_0087_, w_0342_, w_0777_);
not (w_0628_, in2[1]);
or (w_0333_, w_0527_, w_0793_);
and (w_0328_, w_0030_, w_0008_);
or (w_0035_, w_0839_, w_0767_);
and (w_0550_, w_0466_, w_0566_);
and (out7[1], w_0190_, w_0098_);
or (w_0179_, w_0406_, w_0540_);
and (w_0385_, w_0238_, w_0604_);
not (w_0015_, w_0485_);
or (w_0864_, w_0284_, w_0745_);
and (w_0792_, w_0000_, w_0667_);
and (w_0124_, w_0750_, w_0507_);
and (w_0051_, w_0073_, w_0081_);
and (w_0767_, w_0256_, w_0090_);
and (w_0488_, w_0595_, w_0714_);
or (w_0472_, w_0694_, out12[0]);
or (w_0408_, in6[1], in7[1]);
or (w_0508_, w_0103_, w_0395_);
and (w_0576_, w_0750_, w_0633_);
and (w_0849_, in6[2], in7[2]);
not (w_0209_, w_0081_);
and (w_0242_, w_0299_, w_0258_);
and (w_0327_, w_0661_, w_0108_);
not (w_0774_, w_0110_);
not (w_0784_, in8[0]);
or (w_0595_, w_0354_, w_0601_);
and (w_0225_, w_0192_, w_0127_);
and (w_0039_, w_0297_, w_0494_);
and (w_0460_, w_0067_, w_0810_);
and (w_0666_, w_0687_, w_0706_);
and (w_0808_, w_0085_, w_0560_);
or (w_0598_, w_0861_, w_0556_);
and (w_0645_, w_0405_, w_0296_);
and (w_0497_, w_0338_, w_0378_);
and (w_0625_, w_0486_, w_0532_);
not (w_0384_, in13[3]);
or (w_0768_, w_0375_, w_0700_);
and (w_0147_, in8[2], in9[2]);
or (out12[0], w_0540_, w_0460_);
or (w_0193_, w_0594_, w_0592_);
and (w_0501_, w_0861_, w_0556_);
or (w_0127_, in8[3], in9[3]);
or (w_0083_, w_0188_, w_0707_);
not (w_0106_, w_0856_);
and (w_0827_, w_0854_, w_0101_);
or (out10[1], w_0690_, w_0573_);
or (w_0072_, w_0352_, w_0331_);
not (w_0305_, w_0846_);
and (w_0105_, w_0103_, w_0531_);
not (w_0049_, w_0250_);
not (w_0803_, in6[2]);
not (w_0503_, w_0020_);
or (w_0043_, w_0006_, w_0661_);
not (w_0524_, w_0707_);
or (w_0091_, w_0838_, w_0206_);
not (w_0824_, in4[2]);
not (w_0025_, w_0121_);
and (w_0189_, w_0813_, w_0650_);
or (w_0151_, w_0412_, w_0154_);
and (w_0532_, w_0845_, w_0580_);
not (w_0080_, w_0164_);
and (w_0704_, w_0284_, w_0745_);
or (w_0236_, w_0327_, w_0644_);
or (w_0182_, w_0302_, w_0800_);
and (w_0115_, w_0461_, w_0697_);
not (w_0685_, w_0792_);
and (w_0291_, w_0815_, w_0010_);
or (w_0850_, in11[0], in12[0]);
or (w_0070_, in5[2], w_0723_);
or (w_0420_, w_0306_, w_0191_);
and (w_0137_, w_0153_, w_0194_);
and (w_0082_, w_0170_, w_0359_);
or (w_0279_, w_0362_, w_0757_);
and (w_0536_, in6[1], in7[1]);
or (w_0266_, w_0661_, w_0108_);
or (w_0424_, w_0691_, w_0227_);
or (w_0626_, in11[1], in12[1]);
or (out9[1], w_0164_, w_0385_);
not (w_0778_, w_0108_);
or (w_0559_, w_0771_, w_0561_);
or (w_0796_, w_0776_, w_0360_);
and (w_0037_, in4[0], w_0114_);
or (w_0350_, w_0290_, w_0544_);
or (w_0668_, in3[2], w_0189_);
or (w_0119_, w_0506_, w_0325_);
not (w_0830_, in11[0]);
or (w_0058_, w_0389_, w_0781_);
or (w_0798_, in8[2], in9[2]);
and (w_0199_, in13[3], w_0521_);
or (w_0251_, w_0297_, w_0058_);
or (w_0600_, w_0200_, w_0274_);
and (w_0691_, w_0834_, w_0383_);
or (w_0800_, w_0348_, w_0169_);
or (w_0548_, w_0084_, w_0330_);
and (w_0028_, w_0481_, w_0559_);
or (w_0330_, w_0337_, w_0458_);
or (out12[3], w_0454_, w_0051_);
or (w_0483_, w_0265_, w_0666_);
or (w_0036_, w_0476_, w_0762_);
not (w_0309_, w_0063_);
not (w_0776_, in13[1]);
or (w_0276_, w_0399_, w_0320_);
and (w_0614_, w_0097_, w_0603_);
and (w_0777_, w_0165_, w_0474_);
and (w_0195_, w_0638_, w_0220_);
and (w_0323_, w_0178_, w_0172_);
or (w_0138_, w_0102_, w_0373_);
or (w_0572_, w_0338_, w_0378_);
or (w_0398_, w_0731_, w_0817_);
or (w_0660_, w_0016_, w_0432_);
and (w_0842_, w_0333_, w_0841_);
and (w_0107_, w_0343_, w_0615_);
or (w_0571_, w_0386_, w_0124_);
or (w_0526_, w_0339_, w_0715_);
and (w_0673_, w_0432_, w_0073_);
and (w_0586_, w_0168_, w_0712_);
and (w_0793_, w_0367_, w_0434_);
not (w_0504_, w_0072_);
and (w_0678_, w_0581_, w_0093_);
and (w_0461_, w_0251_, w_0864_);
or (w_0823_, w_0209_, w_0235_);
or (out9[2], w_0425_, w_0624_);
or (w_0014_, w_0131_, w_0821_);
or (w_0553_, w_0536_, w_0126_);
or (out2[0], w_0608_, w_0843_);
not (w_0126_, w_0408_);
or (w_0763_, in10[2], w_0790_);
or (w_0387_, w_0758_, w_0071_);
not (w_0506_, in10[0]);
or (w_0097_, w_0546_, w_0361_);
and (w_0237_, w_0302_, w_0446_);
and (w_0156_, out8[1], w_0401_);
or (w_0254_, w_0131_, w_0029_);
or (out6[0], w_0181_, w_0047_);
or (w_0042_, w_0233_, w_0267_);
or (w_0670_, w_0298_, w_0565_);
or (w_0250_, in10[0], w_0682_);
and (w_0566_, w_0688_, w_0078_);
or (w_0136_, w_0851_, w_0357_);
not (w_0733_, in6[0]);
or (out2[1], w_0779_, w_0567_);
and (w_0362_, w_0100_, w_0121_);
and (w_0636_, in10[3], w_0605_);
not (w_0176_, w_0667_);
and (w_0314_, w_0119_, w_0468_);
not (w_0574_, w_0071_);
and (w_0381_, w_0595_, w_0060_);
or (w_0771_, w_0112_, w_0142_);
or (w_0810_, w_0406_, w_0645_);
not (w_0740_, w_0090_);
and (w_0432_, w_0538_, w_0436_);
and (w_0677_, w_0754_, w_0643_);
and (w_0465_, w_0663_, w_0616_);
not (w_0372_, in8[1]);
not (w_0310_, w_0143_);
not (w_0396_, w_0114_);
or (w_0841_, w_0275_, w_0558_);
and (w_0514_, w_0761_, w_0526_);
or (out12[2], w_0322_, w_0451_);
and (w_0535_, w_0545_, w_0074_);
or (w_0365_, out8[2], w_0156_);
or (w_0786_, w_0179_, w_0271_);
not (w_0450_, w_0318_);
and (w_0317_, w_0452_, w_0031_);
not (w_0659_, w_0763_);
and (w_0268_, w_0241_, w_0719_);
not (w_0402_, w_0100_);
and (w_0593_, w_0386_, w_0124_);
or (w_0414_, w_0824_, w_0635_);
or (w_0580_, in5[0], w_0318_);
not (w_0382_, w_0664_);
and (w_0130_, in1[2], in2[2]);
and (w_0271_, w_0007_, w_0587_);
not (w_0040_, in10[1]);
or (w_0557_, in14[1], w_0435_);
and (w_0644_, w_0027_, w_0198_);
and (w_0486_, w_0765_, w_0260_);
not (w_0223_, w_0606_);
and (w_0419_, in11[3], in12[3]);
or (w_0719_, w_0452_, w_0535_);
not (w_0411_, w_0013_);
or (w_0431_, w_0111_, w_0221_);
not (w_0590_, w_0172_);
or (w_0215_, w_0570_, w_0444_);
not (w_0229_, w_0681_);
or (w_0835_, w_0288_, w_0116_);
and (w_0710_, in1[0], w_0691_);
or (w_0795_, w_0780_, w_0056_);
or (w_0654_, w_0550_, w_0797_);
or (w_0094_, w_0345_, w_0278_);
or (w_0163_, w_0207_, w_0609_);
and (w_0388_, in6[0], in7[0]);
or (w_0603_, w_0467_, w_0456_);
not (w_0085_, w_0131_);
not (w_0141_, in13[0]);
not (w_0657_, w_0426_);
or (w_0485_, w_0006_, w_0694_);
or (w_0122_, w_0689_, w_0649_);
or (w_0102_, w_0175_, w_0376_);
or (w_0753_, w_0311_, w_0739_);
and (w_0783_, w_0643_, w_0183_);
not (w_0056_, w_0028_);
not (w_0245_, w_0602_);
or (w_0173_, w_0453_, w_0150_);
and (w_0689_, w_0157_, w_0254_);
and (w_0265_, in11[1], in12[1]);
or (w_0718_, w_0483_, w_0347_);
not (w_0500_, w_0561_);
or (w_0358_, w_0789_, w_0829_);
or (w_0481_, w_0086_, w_0500_);
not (w_0709_, w_0332_);
and (w_0794_, w_0621_, w_0164_);
or (w_0027_, w_0825_, w_0094_);
and (w_0118_, in5[2], w_0723_);
and (w_0348_, in13[1], w_0057_);
not (w_0160_, w_0200_);
or (w_0413_, w_0795_, w_0279_);
not (w_0534_, w_0670_);
and (w_0620_, w_0748_, w_0513_);
and (w_0084_, w_0119_, w_0250_);
or (w_0120_, w_0576_, w_0574_);
or (w_0546_, w_0784_, w_0300_);
and (w_0779_, w_0377_, w_0358_);
or (w_0201_, w_0055_, w_0484_);
not (w_0165_, w_0130_);
not (w_0817_, w_0683_);
and (w_0711_, w_0365_, w_0400_);
and (out7[0], w_0647_, w_0457_);
and (w_0764_, w_0859_, w_0309_);
not (w_0479_, w_0647_);
or (w_0101_, in6[2], in7[2]);
and (w_0298_, in8[1], in9[1]);
not (w_0363_, w_0105_);
and (w_0181_, w_0480_, w_0209_);
or (w_0100_, w_0130_, w_0087_);
and (w_0428_, w_0795_, w_0279_);
and (w_0748_, w_0662_, w_0493_);
and (w_0702_, w_0805_, w_0548_);
and (w_0034_, w_0000_, w_0405_);
not (w_0729_, in10[2]);
and (w_0099_, w_0042_, w_0786_);
not (w_0721_, in12[0]);
or (w_0617_, w_0820_, w_0462_);
and (w_0676_, w_0754_, w_0184_);
or (w_0627_, w_0453_, w_0698_);
or (out4[0], w_0242_, w_0498_);
or (w_0155_, w_0699_, w_0015_);
and (w_0286_, in14[0], w_0237_);
and (w_0487_, w_0022_, w_0703_);
not (w_0492_, w_0668_);
or (w_0074_, w_0391_, w_0743_);
and (w_0739_, w_0215_, w_0511_);
or (w_0180_, w_0631_, w_0551_);
not (w_0696_, w_0398_);
or (w_0637_, w_0064_, w_0021_);
not (w_0186_, w_0017_);
not (w_0148_, w_0453_);
and (w_0567_, w_0738_, w_0392_);
not (w_0032_, w_0167_);
not (w_0541_, w_0070_);
and (w_0613_, w_0671_, w_0545_);
and (w_0061_, w_0045_, w_0425_);
and (w_0543_, w_0648_, w_0716_);
or (w_0243_, w_0669_, w_0277_);
or (w_0041_, w_0037_, w_0554_);
or (w_0805_, w_0273_, w_0437_);
and (w_0860_, w_0759_, w_0408_);
or (w_0692_, w_0145_, w_0282_);
or (w_0641_, w_0727_, w_0336_);
and (w_0862_, w_0494_, w_0011_);
not (w_0132_, w_0078_);
and (w_0573_, in1[1], w_0058_);
or (w_0001_, w_0433_, w_0355_);
or (w_0296_, w_0376_, w_0223_);
and (w_0467_, in8[0], in9[0]);
or (w_0129_, w_0391_, w_0482_);
or (w_0569_, w_0215_, w_0511_);
or (w_0499_, w_0118_, w_0509_);
and (w_0158_, w_0483_, w_0347_);
and (w_0112_, in4[2], w_0678_);
not (w_0221_, w_0470_);
not (w_0315_, w_0278_);
and (w_0207_, w_0854_, w_0091_);
and (w_0240_, w_0218_, w_0418_);
and (w_0444_, w_0288_, w_0116_);
or (w_0701_, w_0748_, w_0513_);
and (w_0683_, w_0110_, w_0660_);
or (w_0185_, w_0199_, w_0370_);
not (w_0178_, w_0053_);
or (w_0312_, w_0791_, w_0623_);
or (w_0020_, w_0199_, w_0319_);
and (w_0621_, w_0201_, w_0247_);
or (w_0104_, in8[0], in9[0]);
or (w_0244_, w_0245_, w_0162_);
or (w_0410_, w_0112_, w_0106_);
and (w_0162_, w_0747_, w_0799_);
and (w_0511_, w_0415_, w_0763_);
or (w_0334_, w_0089_, w_0768_);
or (w_0520_, w_0186_, w_0503_);
and (w_0339_, w_0091_, w_0146_);
or (w_0293_, in8[1], in9[1]);
or (out1[0], w_0785_, w_0632_);
and (w_0169_, w_0776_, w_0360_);
or (w_0684_, w_0490_, w_0423_);
not (w_0459_, in9[1]);
and (w_0561_, w_0059_, w_0448_);
not (w_0383_, w_0781_);
and (w_0456_, w_0826_, w_0293_);
and (w_0406_, w_0220_, w_0441_);
or (w_0329_, w_0836_, w_0770_);
or (w_0671_, w_0125_, w_0728_);
and (w_0303_, w_0692_, w_0280_);
or (w_0466_, w_0111_, w_0158_);
or (w_0184_, in3[1], w_0674_);
not (w_0772_, w_0260_);
or (w_0661_, w_0563_, w_0246_);
or (w_0121_, w_0249_, w_0326_);
and (w_0052_, w_0381_, w_0155_);
or (w_0211_, w_0365_, w_0400_);
or (out7[2], w_0262_, w_0079_);
not (w_0395_, w_0442_);
or (w_0741_, w_0687_, w_0706_);
not (w_0024_, w_0294_);
or (w_0059_, w_0402_, w_0025_);
or (w_0502_, w_0173_, w_0522_);
and (w_0249_, in3[2], w_0189_);
and (w_0652_, w_0658_, w_0542_);
not (w_0135_, w_0240_);
not (w_0609_, w_0734_);
and (w_0089_, w_0630_, w_0439_);
or (w_0359_, w_0816_, w_0487_);
or (w_0369_, w_0426_, w_0477_);
or (w_0662_, w_0367_, w_0434_);
or (w_0427_, w_0018_, w_0272_);
and (w_0435_, w_0182_, w_0196_);
not (w_0021_, w_0397_);
and (w_0002_, w_0176_, w_0252_);
and (w_0554_, w_0329_, w_0088_);
not (w_0843_, w_0510_);
and (w_0623_, w_0680_, w_0751_);
and (w_0131_, w_0480_, w_0137_);
and (w_0563_, w_0084_, w_0330_);
or (w_0801_, w_0203_, w_0656_);
and (w_0069_, w_0694_, out12[0]);
or (w_0425_, w_0465_, w_0248_);
and (w_0743_, w_0671_, w_0397_);
not (w_0228_, w_0837_);
not (w_0308_, w_0810_);
not (w_0757_, w_0481_);
not (w_0829_, w_0236_);
and (w_0476_, in1[1], w_0715_);
or (w_0747_, w_0496_, w_0205_);
or (w_0422_, w_0611_, w_0013_);
not (w_0728_, w_0204_);
or (out5[0], w_0381_, w_0525_);
or (w_0183_, w_0077_, w_0676_);
or (w_0170_, w_0478_, w_0185_);
or (w_0149_, w_0118_, w_0541_);
or (w_0418_, in14[0], w_0237_);
and (w_0527_, w_0036_, w_0128_);
not (w_0855_, w_0617_);
or (w_0579_, w_0029_, w_0693_);
not (w_0144_, in14[1]);
and (w_0594_, w_0166_, w_0471_);
and (w_0140_, w_0802_, w_0096_);
and (w_0610_, w_0773_, w_0668_);
or (w_0630_, w_0144_, w_0575_);
or (w_0022_, w_0384_, w_0654_);
or (w_0469_, w_0134_, w_0403_);
or (w_0717_, w_0593_, w_0695_);
and (w_0638_, w_0520_, w_0120_);
not (w_0599_, w_0224_);
not (w_0306_, in11[2]);
or (w_0171_, w_0722_, w_0304_);
not (w_0054_, w_0012_);
not (w_0744_, w_0210_);
and (w_0370_, w_0384_, w_0654_);
or (w_0340_, w_0640_, w_0562_);
or (w_0720_, in10[3], w_0605_);
or (out9[0], w_0073_, w_0081_);
or (w_0675_, w_0327_, w_0393_);
and (w_0782_, w_0339_, w_0129_);
not (w_0331_, w_0138_);
not (w_0076_, out8[1]);
or (w_0342_, w_0187_, w_0066_);
or (w_0646_, in1[2], w_0734_);
or (out1[1], w_0069_, w_0019_);
and (out11[2], w_0193_, w_0211_);
and (w_0787_, in14[2], w_0784_);
or (w_0198_, w_0016_, w_0299_);
and (w_0341_, w_0380_, w_0858_);
and (w_0715_, w_0809_, w_0243_);
and (w_0693_, w_0672_, w_0014_);
or (w_0371_, w_0351_, w_0063_);
or (w_0390_, w_0665_, w_0107_);
not (w_0393_, w_0266_);
not (w_0214_, w_0626_);
and (w_0203_, w_0796_, w_0182_);
or (w_0856_, in4[2], w_0678_);
and (w_0528_, w_0173_, w_0522_);
and (w_0033_, w_0388_, w_0860_);
and (w_0785_, w_0631_, w_0551_);
and (w_0591_, w_0629_, w_0627_);
or (w_0615_, in1[0], w_0480_);
and (w_0407_, w_0203_, w_0656_);
not (w_0192_, w_0611_);
not (w_0445_, in5[0]);
not (w_0290_, in14[2]);
or (out6[2], w_0862_, w_0061_);
or (w_0259_, w_0702_, w_0778_);
not (w_0447_, w_0806_);
or (w_0857_, w_0461_, w_0697_);
and (w_0368_, in1[2], w_0734_);
and (w_0285_, w_0801_, w_0598_);
and (w_0513_, w_0424_, w_0255_);
and (w_0294_, w_0653_, w_0190_);
or (w_0745_, w_0710_, w_0755_);
and (w_0714_, w_0469_, w_0229_);
not (w_0780_, w_0499_);
and (w_0275_, w_0058_, w_0244_);
and (w_0263_, w_0290_, in8[0]);
or (w_0010_, in1[1], w_0253_);
or (out6[1], w_0847_, w_0794_);
or (w_0397_, in5[1], w_0204_);
or (w_0026_, w_0497_, w_0428_);
or (w_0438_, w_0625_, w_0268_);
and (w_0790_, w_0517_, w_0732_);
not (w_0191_, in12[2]);
not (w_0746_, w_0412_);
or (w_0575_, w_0324_, w_0832_);
or (w_0177_, in13[1], w_0057_);
or (w_0161_, w_0139_, w_0374_);
and (w_0451_, w_0714_, w_0694_);
or (w_0012_, w_0339_, w_0129_);
and (w_0570_, in10[1], w_0614_);
and (w_0366_, w_0006_, w_0661_);
not (w_0353_, w_0799_);
or (w_0316_, in1[2], w_0494_);
not (w_0019_, w_0472_);
and (w_0663_, w_0413_, w_0572_);
not (w_0048_, w_0699_);
or (w_0650_, w_0342_, w_0777_);
or (w_0016_, w_0034_, w_0195_);
and (w_0453_, w_0432_, w_0494_);
not (w_0218_, w_0286_);
or (w_0592_, w_0512_, w_0588_);
or (w_0234_, w_0516_, w_0363_);
not (w_0616_, w_0766_);
not (w_0374_, w_0643_);
and (out3[0], w_0823_, w_0749_);
and (w_0781_, w_0046_, w_0535_);
and (w_0073_, w_0455_, w_0568_);
or (w_0581_, w_0677_, w_0597_);
not (w_0233_, w_0179_);
or (w_0302_, w_0141_, w_0744_);
not (w_0416_, in7[1]);
and (w_0723_, w_0050_, w_0151_);
not (w_0235_, w_0579_);
or (w_0196_, w_0430_, w_0113_);
not (w_0389_, w_0834_);
or (w_0474_, in1[2], in2[2]);
and (w_0347_, w_0420_, w_0470_);
not (w_0680_, in14[3]);
and (w_0326_, w_0161_, w_0610_);
or (w_0577_, in1[1], in2[1]);
not (w_0241_, w_0188_);
or (w_0386_, w_0375_, w_0352_);
and (w_0769_, w_0144_, w_0575_);
not (w_0454_, out9[0]);
and (w_0762_, w_0018_, w_0272_);
or (w_0669_, w_0064_, w_0863_);
or (w_0596_, in3[0], w_0105_);
and (w_0515_, w_0630_, w_0557_);
and (w_0821_, w_0323_, w_0595_);
or (w_0597_, w_0249_, w_0492_);
and (w_0168_, w_0415_, w_0713_);
and (w_0164_, w_0109_, w_0600_);
or (w_0457_, w_0137_, w_0099_);
not (w_0145_, in11[1]);
not (w_0345_, w_0281_);
and (w_0288_, in10[0], w_0682_);
and (w_0391_, in5[0], w_0318_);
or (w_0518_, w_0736_, w_0143_);
and (w_0811_, in4[1], w_0783_);
or (w_0612_, w_0046_, w_0734_);
not (w_0005_, w_0714_);
not (w_0491_, in1[2]);
and (w_0484_, w_0032_, w_0519_);
and (w_0373_, w_0350_, w_0814_);
not (w_0853_, w_0627_);
or (w_0000_, w_0364_, w_0337_);
or (w_0686_, w_0084_, w_0240_);
or (w_0647_, w_0595_, w_0258_);
not (w_0822_, w_0782_);
and (w_0154_, w_0414_, w_0856_);
not (w_0289_, w_0320_);
not (w_0516_, in3[0]);
or (w_0732_, w_0670_, w_0224_);
and (w_0766_, w_0163_, w_0109_);
and (w_0003_, w_0837_, w_0679_);
and (w_0558_, w_0691_, w_0227_);
and (w_0690_, w_0727_, w_0691_);
not (w_0820_, w_0083_);
or (w_0280_, w_0380_, w_0858_);
and (w_0167_, w_0753_, w_0475_);
or (w_0090_, w_0747_, w_0799_);
or (w_0602_, w_0491_, w_0045_);
not (w_0417_, w_0646_);
not (w_0463_, w_0274_);
or (w_0665_, w_0774_, w_0696_);
and (w_0045_, w_0822_, w_0012_);
or (w_0533_, w_0388_, w_0772_);
or (w_0664_, in10[1], w_0614_);
or (w_0255_, w_0058_, w_0244_);
and (w_0509_, w_0669_, w_0277_);
or (w_0470_, in11[2], in12[2]);
and (w_0224_, w_0001_, w_0798_);
not (w_0565_, w_0097_);
and (w_0863_, w_0391_, w_0743_);
or (w_0587_, w_0806_, w_0504_);
and (w_0505_, w_0137_, w_0005_);
not (w_0038_, w_0107_);
or (w_0252_, w_0422_, w_0607_);
or (w_0197_, w_0714_, w_0694_);
not (w_0458_, w_0387_);
or (w_0044_, w_0638_, w_0220_);
not (w_0640_, w_0343_);
or (w_0584_, w_0228_, w_0673_);
not (w_0295_, w_0720_);
and (w_0062_, w_0208_, w_0270_);
or (w_0585_, w_0147_, w_0844_);
or (w_0446_, in13[0], w_0210_);
and (w_0552_, w_0864_, w_0502_);
and (w_0838_, w_0759_, w_0828_);
not (w_0844_, w_0517_);
and (w_0053_, w_0806_, w_0533_);
and (w_0496_, in1[1], w_0253_);
or (w_0292_, w_0017_, w_0020_);
or (w_0839_, w_0762_, w_0115_);
or (w_0523_, w_0065_, w_0789_);
or (w_0845_, w_0445_, w_0450_);
not (w_0727_, in1[1]);
and (w_0057_, w_0280_, w_0741_);
not (w_0736_, w_0589_);
not (w_0455_, w_0578_);
and (w_0299_, w_0281_, w_0315_);
and (w_0755_, w_0297_, w_0058_);
and (w_0522_, w_0251_, w_0301_);
or (w_0212_, w_0321_, w_0307_);
not (w_0760_, w_0313_);
and (w_0649_, w_0369_, w_0808_);
and (w_0134_, w_0007_, w_0042_);
or (w_0281_, in14[3], in8[1]);
or (w_0854_, w_0803_, w_0222_);
and (w_0512_, w_0839_, w_0767_);
and (w_0274_, w_0163_, w_0612_);
or (w_0468_, w_0570_, w_0382_);
and (w_0332_, w_0437_, w_0002_);
or (w_0480_, w_0053_, w_0590_);
or (w_0108_, w_0787_, w_0263_);
not (w_0688_, w_0419_);
and (w_0174_, w_0159_, w_0390_);
and (w_0583_, w_0722_, w_0304_);
or (w_0109_, w_0160_, w_0463_);
and (w_0478_, w_0171_, w_0801_);
or (w_0448_, w_0100_, w_0121_);
and (w_0248_, w_0026_, w_0766_);
and (w_0364_, w_0017_, w_0020_);
not (w_0840_, in3[1]);
and (out11[1], w_0471_, w_0547_);
or (w_0304_, w_0158_, w_0213_);
and (w_0337_, w_0758_, w_0071_);
and (w_0440_, w_0582_, w_0827_);
and (w_0629_, w_0657_, w_0429_);
or (w_0815_, w_0727_, w_0621_);
and (w_0437_, w_0120_, w_0387_);
and (w_0716_, w_0685_, w_0555_);
and (w_0150_, w_0075_, w_0853_);
and (w_0143_, in7[1], in2[1]);
or (w_0321_, w_0529_, w_0396_);
and (w_0377_, w_0731_, w_0043_);
and (w_0220_, w_0542_, w_0835_);
and (w_0611_, in8[3], in9[3]);
and (w_0376_, w_0286_, w_0515_);
and (w_0799_, w_0602_, w_0316_);
and (w_0064_, in5[1], w_0204_);
and (w_0324_, w_0430_, w_0113_);
or (w_0093_, w_0161_, w_0610_);
and (w_0378_, w_0059_, w_0481_);
or (w_0394_, w_0150_, w_0591_);
not (w_0462_, w_0514_);
or (w_0346_, w_0409_, w_0231_);
or (w_0449_, w_0162_, w_0740_);
or (w_0861_, w_0348_, w_0324_);
and (w_0707_, w_0625_, w_0268_);
or (w_0738_, w_0366_, w_0622_);
or (w_0837_, w_0432_, w_0073_);
or (w_0538_, in7[2], in2[2]);
and (w_0065_, w_0016_, w_0299_);
not (w_0357_, w_0469_);
not (w_0529_, in4[0]);
not (w_0261_, w_0823_);
not (w_0355_, in9[2]);
or (w_0172_, w_0806_, w_0533_);
or (w_0301_, in1[0], w_0691_);
not (w_0731_, w_0366_);
and (w_0825_, w_0044_, w_0833_);
or (w_0405_, w_0444_, w_0314_);
or (w_0735_, w_0006_, w_0714_);
or (w_0544_, w_0501_, w_0407_);
or (w_0604_, w_0648_, w_0716_);
or (w_0712_, w_0636_, w_0295_);
and (w_0601_, in7[0], in2[0]);
and (w_0674_, w_0508_, w_0335_);
or (w_0742_, w_0099_, w_0631_);
and (w_0651_, w_0857_, w_0427_);
and (w_0319_, w_0816_, w_0487_);
or (w_0582_, w_0536_, w_0033_);
or (out10[2], w_0464_, w_0092_);
or (w_0606_, w_0286_, w_0515_);
or (w_0159_, w_0257_, w_0038_);
or (w_0287_, w_0499_, w_0028_);
and (w_0313_, w_0653_, w_0735_);
not (w_0761_, w_0489_);
or (w_0751_, w_0319_, w_0217_);
and (w_0204_, w_0212_, w_0041_);
or (out10[0], w_0039_, w_0804_);
not (w_0635_, w_0678_);
not (w_0482_, w_0580_);
and (w_0320_, w_0009_, w_0291_);
not (w_0622_, w_0043_);
and (w_0116_, w_0658_, w_0664_);
or (w_0231_, w_0419_, w_0132_);
or (out3[1], w_0812_, w_0756_);
or (w_0360_, w_0666_, w_0341_);
not (w_0194_, w_0601_);
or (w_0380_, w_0830_, w_0721_);
and (w_0246_, w_0273_, w_0437_);
and (w_0079_, w_0294_, w_0003_);
and (w_0029_, w_0523_, w_0216_);
and (w_0352_, w_0102_, w_0373_);
and (w_0175_, in14[1], w_0435_);
not (w_0349_, w_0636_);
or (w_0128_, w_0417_, w_0368_);
not (w_0267_, w_0271_);
and (w_0642_, w_0709_, w_0404_);
or (w_0834_, w_0046_, w_0535_);
or (w_0166_, w_0552_, w_0708_);
not (w_0404_, w_0619_);
or (w_0078_, in11[3], in12[3]);
and (out11[0], w_0076_, w_0655_);
or (w_0631_, w_0625_, w_0473_);
or (w_0759_, w_0775_, w_0416_);
and (w_0113_, w_0796_, w_0177_);
and (w_0734_, w_0795_, w_0287_);
and (w_0789_, w_0327_, w_0644_);
and (w_0096_, w_0048_, w_0485_);
or (w_0658_, w_0040_, w_0239_);
or (w_0542_, w_0119_, w_0468_);
not (w_0361_, w_0456_);
not (w_0095_, in2[0]);
not (w_0775_, in6[1]);
and (w_0077_, in3[0], w_0105_);
or (w_0726_, w_0083_, w_0514_);
not (w_0773_, w_0249_);
and (w_0797_, w_0409_, w_0231_);
or (w_0858_, w_0265_, w_0214_);
and (w_0071_, w_0520_, w_0292_);
or (w_0256_, w_0530_, w_0353_);
or (w_0788_, w_0009_, w_0291_);
and (w_0852_, w_0825_, w_0094_);
and (w_0272_, w_0641_, w_0846_);
not (w_0232_, w_0676_);
or (w_0517_, w_0534_, w_0599_);
and (w_0092_, w_0491_, w_0715_);
and (w_0549_, w_0398_, w_0564_);
not (w_0060_, w_0631_);
not (w_0239_, w_0614_);
and (w_0477_, w_0518_, w_0621_);
not (w_0157_, w_0369_);
or (w_0826_, w_0372_, w_0459_);
or (w_0202_, w_0311_, w_0659_);
or (w_0750_, w_0680_, w_0751_);
and (w_0152_, w_0350_, w_0334_);
and (w_0006_, w_0589_, w_0310_);
and (w_0540_, w_0133_, w_0308_);
and (w_0737_, w_0037_, w_0554_);
and (w_0672_, w_0027_, w_0023_);
or (w_0814_, in14[2], w_0285_);
or (w_0846_, in1[1], w_0715_);
not (w_0530_, w_0747_);
and (w_0318_, w_0321_, w_0123_);
and (w_0806_, w_0713_, w_0569_);
or (w_0031_, w_0167_, w_0586_);
or (w_0023_, w_0259_, w_0264_);
and (w_0699_, w_0006_, w_0694_);
not (w_0848_, w_0790_);
or (w_0050_, w_0746_, w_0410_);
or (w_0098_, w_0479_, w_0313_);
and (w_0311_, in10[2], w_0790_);
not (w_0730_, w_0368_);
and (w_0111_, in11[2], in12[2]);
and (w_0578_, w_0136_, w_0642_);
or (w_0634_, out8[2], w_0269_);
not (w_0257_, w_0665_);
or (out5[1], w_0140_, w_0052_);
or (w_0507_, in14[3], w_0082_);
not (w_0813_, w_0087_);
or (w_0403_, w_0851_, w_0068_);
not (w_0421_, w_0101_);
or (w_0531_, in1[0], in2[0]);
and (w_0556_, w_0171_, w_0283_);
not (w_0238_, w_0543_);
not (w_0300_, in9[0]);
not (w_0297_, in1[0]);
or (w_0007_, w_0447_, w_0072_);
and (w_0752_, in1[0], in2[0]);
or (w_0103_, w_0297_, w_0095_);
or (w_0749_, w_0081_, w_0579_);
and (w_0068_, w_0031_, w_0717_);
and (w_0562_, w_0665_, w_0107_);
and (w_0791_, in14[3], w_0082_);
and (w_0401_, w_0166_, w_0004_);
not (w_0322_, w_0197_);
or (w_0819_, w_0258_, w_0060_);
and (w_0804_, in1[0], w_0045_);
or (w_0260_, in6[0], in7[0]);
and (w_0081_, w_0617_, w_0726_);
and (w_0681_, w_0134_, w_0403_);
and (w_0832_, w_0302_, w_0800_);
or (w_0379_, w_0175_, w_0769_);
and (w_0205_, w_0340_, w_0010_);
not (w_0133_, w_0067_);
not (w_0490_, w_0538_);
or (w_0190_, w_0647_, w_0760_);
or (w_0017_, w_0419_, w_0550_);
or (w_0146_, w_0582_, w_0827_);
and (w_0618_, w_0055_, w_0484_);
not (w_0433_, in8[2]);
and (w_0230_, w_0765_, w_0553_);
or (w_0807_, w_0727_, w_0628_);
not (w_0770_, w_0783_);
or (w_0859_, w_0164_, w_0122_);
and (w_0434_, w_0646_, w_0730_);
and (w_0210_, w_0380_, w_0850_);
not (w_0679_, w_0673_);
and (w_0687_, in11[0], in12[0]);
and (w_0047_, w_0323_, w_0081_);
or (w_0088_, in4[1], w_0783_);
or (w_0697_, w_0476_, w_0305_);
and (w_0423_, in7[2], in2[2]);
and (w_0498_, w_0094_, w_0099_);
and (w_0851_, w_0484_, w_0724_);
not (w_0836_, in4[1]);
or (w_0117_, w_0585_, w_0225_);
not (w_0338_, w_0795_);
or (w_0439_, w_0218_, w_0379_);
or (w_0200_, w_0489_, w_0855_);
or (w_0429_, w_0369_, w_0808_);
or (w_0335_, w_0752_, w_0442_);
and (w_0605_, w_0411_, w_0117_);
or (w_0273_, w_0288_, w_0049_);
and (w_0682_, w_0546_, w_0104_);
and (w_0708_, w_0788_, w_0289_);
or (w_0653_, w_0518_, w_0005_);
and (w_0847_, w_0253_, w_0080_);
not (w_0356_, in7[0]);
or (out4[1], w_0505_, w_0488_);
and (w_0756_, w_0823_, w_0764_);
or (w_0560_, w_0672_, w_0014_);
not (w_0125_, in5[1]);
or (w_0555_, w_0000_, w_0667_);
and (w_0473_, w_0533_, w_0129_);
or (w_0153_, in7[0], in2[0]);
or (w_0643_, w_0234_, w_0232_);
and (w_0262_, w_0024_, w_0584_);
and (w_0269_, w_0552_, w_0708_);
or (w_0030_, w_0842_, w_0620_);
not (w_0336_, w_0715_);
or (w_0816_, w_0219_, w_0501_);
and (w_0430_, in13[0], w_0210_);
not (w_0282_, in12[1]);
and (w_0277_, w_0344_, w_0070_);
and (w_0525_, w_0137_, w_0631_);
not (w_0632_, w_0180_);
and (w_0667_, w_0422_, w_0607_);
not (w_0392_, w_0358_);
and (w_0188_, w_0452_, w_0535_);
or (w_0123_, in4[0], w_0114_);
not (out8[2], w_0166_);
not (w_0086_, w_0771_);
or (w_0828_, w_0765_, w_0553_);
or (w_0545_, w_0845_, w_0637_);
and (w_0551_, w_0067_, w_0686_);
not (w_0258_, w_0099_);
or (w_0206_, w_0849_, w_0421_);
or (w_0270_, w_0512_, w_0711_);
or (w_0493_, w_0036_, w_0128_);
and (w_0227_, w_0602_, w_0256_);
and (w_0442_, w_0807_, w_0577_);
not (w_0722_, in13[2]);
and (out8[0], w_0122_, w_0549_);
or (w_0754_, w_0840_, w_0495_);
not (w_0495_, w_0674_);
and (w_0698_, w_0684_, w_0045_);
not (w_0354_, w_0153_);
and (w_0475_, w_0349_, w_0720_);
or (w_0539_, w_0528_, w_0704_);
not (w_0724_, w_0717_);
or (w_0247_, w_0452_, w_0031_);
and (w_0619_, w_0330_, w_0818_);
not (w_0307_, w_0554_);
not (w_0142_, w_0050_);
and (w_0409_, w_0420_, w_0443_);
or (w_0765_, w_0733_, w_0356_);
or (w_0831_, w_0629_, w_0627_);
or (w_0656_, w_0219_, w_0583_);
and (w_0426_, w_0006_, w_0253_);
or (w_0705_, w_0651_, w_0449_);
or (w_0713_, w_0652_, w_0202_);
or (w_0253_, w_0317_, w_0618_);
and (w_0013_, w_0585_, w_0225_);
endmodule

module sub_module2(
    input wire [1:0] in1,
    input wire [1:0] in2,
    input wire [1:0] in3,
    input wire [1:0] in4,
    input wire [1:0] in5,
    input wire [1:0] in6,
    input wire [1:0] in7,
    input wire [4:0] in8,
    input wire [4:0] in9,
    input wire [4:0] in10,
    input wire [4:0] in11,
    input wire [4:0] in12,
    input wire [4:0] in13,
    input wire [4:0] in14,
    input wire [4:0] in15,
    output wire [1:0] out1,
    output wire [1:0] out2,
    output wire [1:0] out3,
    output wire [1:0] out4,
    output wire [1:0] out5,
    output wire [2:0] out6,
    output wire [2:0] out7,
    output wire [2:0] out8,
    output wire [2:0] out9,
    output wire [2:0] out10,
    output wire [3:0] out11,
    output wire [3:0] out12,
    output wire [3:0] out13,
    output wire [3:0] out14
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
wire w_0945_;
wire w_0946_;
wire w_0947_;
wire w_0948_;
wire w_0949_;
wire w_0950_;
wire w_0951_;
wire w_0952_;
wire w_0953_;
wire w_0954_;
wire w_0955_;
wire w_0956_;
wire w_0957_;
wire w_0958_;
wire w_0959_;
wire w_0960_;
wire w_0961_;
wire w_0962_;
wire w_0963_;
wire w_0964_;
wire w_0965_;
wire w_0966_;
wire w_0967_;
wire w_0968_;
wire w_0969_;
wire w_0970_;
wire w_0971_;
wire w_0972_;
wire w_0973_;
wire w_0974_;
wire w_0975_;
wire w_0976_;
wire w_0977_;
wire w_0978_;
wire w_0979_;
wire w_0980_;
wire w_0981_;
wire w_0982_;
wire w_0983_;
wire w_0984_;
wire w_0985_;
wire w_0986_;
wire w_0987_;
wire w_0988_;
wire w_0989_;
wire w_0990_;
wire w_0991_;
wire w_0992_;
wire w_0993_;
wire w_0994_;
wire w_0995_;
wire w_0996_;
wire w_0997_;
wire w_0998_;
wire w_0999_;
wire w_1000_;
wire w_1001_;
wire w_1002_;
wire w_1003_;
wire w_1004_;
wire w_1005_;
wire w_1006_;
wire w_1007_;
wire w_1008_;
wire w_1009_;
wire w_1010_;
wire w_1011_;
wire w_1012_;
wire w_1013_;
wire w_1014_;
wire w_1015_;
wire w_1016_;
wire w_1017_;
wire w_1018_;
wire w_1019_;
wire w_1020_;
wire w_1021_;
wire w_1022_;
wire w_1023_;
wire w_1024_;
and (w_0703_, w_0593_, w_0012_);
and (w_0011_, w_0477_, w_0810_);
or (w_0644_, w_0217_, w_0567_);
and (w_0173_, w_0459_, w_0479_);
and (w_0744_, w_0856_, w_0717_);
and (w_0392_, w_0700_, w_0198_);
or (w_0522_, w_0844_, w_0483_);
and (w_0681_, in13[1], in12[1]);
or (w_0567_, w_0310_, w_0699_);
and (w_0572_, w_0673_, w_0780_);
not (w_0604_, in9[1]);
and (w_0796_, w_0064_, w_0925_);
and (w_1007_, w_0009_, w_0609_);
and (w_0552_, w_0546_, w_0817_);
and (w_0975_, w_0662_, w_0198_);
and (w_0529_, w_0233_, w_0657_);
and (w_0906_, w_0323_, w_0005_);
and (w_0993_, w_0077_, w_0593_);
or (w_0306_, w_0647_, w_0395_);
or (w_0841_, w_0080_, w_0238_);
and (w_0872_, w_0017_, w_0358_);
and (w_0388_, w_0936_, w_0140_);
or (w_0138_, w_0429_, w_0188_);
and (w_0078_, w_0308_, w_0036_);
or (w_0563_, w_0681_, w_1013_);
or (w_0469_, w_0967_, w_0237_);
or (out8[0], w_0330_, w_0747_);
or (w_0329_, w_0388_, w_0414_);
and (w_0595_, w_0239_, w_0663_);
or (w_0905_, in9[1], in8[1]);
and (w_0556_, w_0315_, w_0046_);
or (w_0320_, w_0111_, w_0671_);
and (w_0311_, w_0650_, w_0299_);
not (w_0083_, w_0723_);
and (w_0150_, w_0501_, w_0923_);
or (w_0626_, w_0034_, w_0267_);
or (w_0615_, in9[4], in8[4]);
and (w_0208_, w_0076_, w_0552_);
and (w_0451_, w_0480_, w_0373_);
or (w_0748_, w_0325_, w_0378_);
or (w_0774_, w_0133_, w_0894_);
not (w_0165_, w_0684_);
or (w_0981_, w_0861_, w_0055_);
and (w_0534_, w_0678_, w_0692_);
and (w_0839_, w_0385_, w_0518_);
or (w_0226_, w_0462_, w_0910_);
not (w_0190_, w_0074_);
and (w_0640_, w_0400_, w_0139_);
and (w_0422_, w_0198_, w_0300_);
and (w_0705_, w_0329_, w_0637_);
or (w_0850_, in15[4], w_0808_);
or (w_0023_, w_0038_, w_1012_);
and (w_1012_, w_0908_, w_0685_);
or (w_0331_, w_0991_, w_0495_);
and (w_0817_, w_0799_, w_0743_);
not (w_0955_, in11[1]);
and (w_0456_, w_0079_, w_0768_);
or (w_0917_, w_0255_, w_0957_);
or (w_0617_, w_0977_, w_0099_);
and (w_0314_, w_0140_, w_0985_);
and (w_1024_, w_0992_, w_0303_);
not (w_0576_, w_0758_);
not (w_0216_, w_0795_);
or (w_0421_, w_0529_, w_0056_);
and (w_0119_, w_0371_, w_0926_);
or (w_0460_, w_0643_, w_0445_);
and (w_0409_, w_0583_, w_0539_);
or (w_0509_, in1[0], in2[0]);
and (w_0056_, w_0737_, w_0770_);
or (w_0006_, w_0828_, w_0963_);
and (w_0585_, w_0326_, w_0783_);
not (w_0713_, w_0289_);
or (w_0740_, in2[0], w_0280_);
or (w_0554_, w_0794_, w_0881_);
and (w_0634_, w_0686_, w_0670_);
or (w_0151_, w_0899_, w_0113_);
and (w_0275_, w_0260_, w_0034_);
and (w_0855_, w_0511_, w_0660_);
or (w_0021_, w_0830_, w_0481_);
and (w_1005_, w_0215_, w_0040_);
or (w_0194_, w_0076_, w_0223_);
or (w_0506_, w_0050_, w_0956_);
not (w_0671_, w_0859_);
or (w_0800_, w_0379_, w_0426_);
and (w_0330_, w_0518_, w_0072_);
and (w_0063_, w_0010_, w_0753_);
not (w_0287_, w_0313_);
and (w_0490_, w_0331_, w_0107_);
not (w_0156_, w_0080_);
not (w_0336_, in11[0]);
or (w_0187_, w_0514_, w_0617_);
or (w_0039_, w_0216_, w_0143_);
not (w_0659_, w_0860_);
and (w_0473_, w_0878_, w_0269_);
or (w_0969_, w_0018_, w_0875_);
and (w_0146_, w_0178_, w_0086_);
and (w_0791_, w_0161_, w_0763_);
not (w_0256_, w_0504_);
or (w_0694_, w_0891_, w_0098_);
and (w_0544_, in10[3], w_1024_);
or (w_0477_, w_0475_, w_0636_);
not (w_1020_, w_0583_);
or (w_0420_, w_0835_, w_0354_);
or (w_0131_, w_0426_, w_0638_);
and (w_0380_, w_0813_, w_0277_);
and (w_0973_, w_0913_, w_0195_);
not (w_1000_, w_1024_);
or (w_0478_, w_0498_, w_0938_);
or (w_0299_, w_0746_, w_0986_);
or (out10[2], w_0380_, w_0573_);
and (w_0164_, w_0111_, w_0341_);
or (w_0048_, w_0090_, w_0759_);
or (w_0847_, w_0656_, w_0304_);
or (w_0300_, w_0338_, w_0053_);
or (w_0553_, w_0083_, w_0121_);
and (w_0862_, w_0547_, w_0904_);
and (w_0831_, w_0746_, w_0986_);
and (w_0565_, w_0813_, w_0362_);
and (w_0970_, in13[0], in12[0]);
not (w_0294_, in15[1]);
or (w_0424_, w_0766_, w_0421_);
or (w_0349_, w_0677_, w_0366_);
or (out3[1], w_0791_, w_0410_);
and (w_0461_, w_0320_, w_0675_);
or (w_0343_, w_0887_, w_0449_);
and (w_0067_, w_0169_, w_0285_);
and (w_0802_, w_0870_, w_0668_);
and (w_0945_, w_0809_, w_0070_);
or (w_0566_, w_0416_, w_0054_);
and (w_0723_, w_0172_, w_0000_);
not (w_0288_, w_0065_);
or (w_0413_, w_0145_, w_0342_);
or (w_0457_, w_0981_, w_0095_);
or (w_0132_, in15[1], w_0634_);
and (w_0837_, w_0187_, w_0168_);
and (w_0716_, w_0404_, w_0161_);
not (w_0394_, w_0136_);
not (w_0536_, w_0490_);
and (w_0260_, w_0784_, w_0485_);
or (w_0933_, w_0017_, w_0737_);
and (w_0951_, w_0821_, w_0591_);
and (w_0784_, w_0312_, w_0441_);
not (w_0211_, w_0446_);
or (w_0755_, w_0997_, w_0028_);
or (w_0890_, w_0724_, w_0311_);
and (w_0961_, in10[4], w_0602_);
or (w_0458_, w_0431_, w_0556_);
and (w_0341_, w_0555_, w_0068_);
or (w_0434_, w_1014_, w_0415_);
and (w_0620_, w_0838_, w_0813_);
and (w_0834_, w_0372_, w_0640_);
and (w_0546_, w_0720_, w_0496_);
or (w_0637_, w_0738_, w_0764_);
or (w_0312_, w_0009_, w_0079_);
or (w_0279_, w_0263_, w_0204_);
not (w_0887_, in14[4]);
and (w_0262_, w_0522_, w_0134_);
or (w_0924_, w_0697_, w_0251_);
and (w_0155_, w_0514_, w_0765_);
or (w_0335_, w_0965_, w_0157_);
and (w_0503_, w_0048_, w_0851_);
and (w_0035_, w_0562_, w_0739_);
and (w_0356_, in9[3], in8[3]);
or (w_0697_, w_0242_, w_0581_);
or (w_0507_, w_0322_, w_0131_);
not (w_0088_, in1[0]);
and (w_0271_, w_0365_, w_0885_);
and (w_0896_, w_0396_, w_0576_);
or (w_0363_, w_1015_, w_0947_);
and (w_0143_, w_0945_, w_0958_);
and (w_0030_, w_0019_, w_0967_);
or (w_0229_, w_0831_, w_0029_);
not (w_0238_, w_0710_);
and (w_0286_, w_0362_, w_0403_);
and (w_0513_, w_0922_, w_0684_);
and (w_0050_, w_0263_, w_0204_);
not (w_0346_, in2[0]);
and (w_0201_, w_0765_, w_0364_);
or (w_0986_, w_0733_, w_1004_);
or (w_0147_, w_0310_, w_0873_);
or (w_0091_, w_0166_, w_0196_);
and (w_0065_, w_0148_, w_0987_);
and (w_0525_, w_0797_, w_0339_);
or (w_0725_, w_0702_, w_0585_);
or (w_0510_, w_0550_, w_0532_);
or (w_0345_, w_0274_, w_0575_);
and (w_0248_, w_0793_, w_0044_);
and (w_0695_, w_0186_, w_0590_);
or (w_0888_, w_0321_, w_0620_);
not (w_0674_, w_0966_);
or (w_0717_, w_0431_, w_0287_);
not (w_0369_, w_0475_);
or (w_0044_, w_0477_, w_0810_);
or (w_0202_, w_0148_, w_0758_);
or (w_0338_, w_0873_, w_0027_);
and (w_0941_, w_0925_, w_0748_);
or (w_0739_, in13[4], in12[4]);
or (w_0234_, w_0243_, w_0757_);
not (w_0564_, w_0628_);
and (w_0956_, w_0170_, w_0007_);
or (w_0932_, w_0716_, w_0253_);
not (w_0500_, in9[3]);
or (w_0470_, w_0177_, w_0228_);
and (w_0533_, w_0343_, w_0624_);
not (w_0562_, w_0687_);
or (w_0570_, w_0945_, w_0274_);
and (w_1016_, w_0159_, w_0026_);
or (w_0465_, w_0857_, w_0823_);
and (w_0222_, w_0723_, w_0229_);
and (w_0383_, w_0932_, w_0682_);
or (w_0389_, w_0673_, w_0161_);
and (w_0535_, w_1001_, w_0997_);
or (out10[0], w_0032_, w_0461_);
or (w_0768_, w_0008_, w_0450_);
or (out1[0], w_0979_, w_0568_);
and (w_0600_, w_0887_, w_0449_);
or (w_0826_, w_0289_, w_0779_);
or (w_0916_, w_0622_, w_0084_);
and (w_0602_, w_0151_, w_0292_);
and (w_0240_, w_0193_, w_0306_);
and (w_0607_, w_0385_, w_0559_);
and (w_0250_, w_0268_, w_0319_);
or (w_0205_, w_0028_, w_1022_);
or (w_0743_, w_0233_, w_0657_);
or (w_0819_, w_0690_, w_0995_);
not (w_0144_, w_0345_);
not (w_0308_, in14[2]);
and (w_0359_, w_0502_, w_0066_);
or (w_0135_, w_0835_, w_1016_);
not (w_0018_, in15[2]);
or (w_0218_, w_0239_, w_0663_);
or (w_0666_, w_0687_, w_0868_);
or (w_0057_, w_1001_, w_0997_);
or (w_0447_, w_0714_, w_0226_);
and (w_0976_, w_0432_, w_1022_);
not (w_0726_, in9[2]);
or (w_0555_, w_0955_, w_0645_);
and (w_0588_, w_0857_, w_0823_);
or (w_0340_, w_0958_, w_0263_);
and (w_0767_, w_0268_, w_0270_);
or (w_0763_, w_0959_, w_0906_);
or (w_0376_, w_0472_, w_0879_);
or (w_0502_, w_0828_, w_1014_);
and (w_0316_, w_0123_, w_0453_);
or (w_0947_, w_0141_, w_0976_);
and (w_0198_, w_0209_, w_0298_);
or (w_0686_, w_0002_, w_0603_);
and (w_0977_, in15[0], w_0824_);
or (out10[1], w_0162_, w_0614_);
or (w_0269_, w_0432_, w_0399_);
and (w_0277_, w_0447_, w_0234_);
or (w_0781_, w_0297_, w_0521_);
and (w_0601_, w_0257_, w_0826_);
and (w_0407_, w_0795_, w_0907_);
and (w_0484_, w_0237_, w_0198_);
and (w_0185_, w_0309_, w_0512_);
or (w_0036_, w_1023_, w_0042_);
and (w_0794_, w_0224_, w_0524_);
and (w_0276_, w_0550_, w_0532_);
and (w_0519_, w_0758_, w_0700_);
and (w_0928_, w_0664_, w_0281_);
or (w_0064_, w_0137_, w_0789_);
not (w_0110_, w_0061_);
or (w_0170_, w_0700_, w_0198_);
and (w_0027_, w_0217_, w_0567_);
and (w_0101_, in14[1], w_0230_);
and (w_0729_, w_0177_, w_0228_);
and (w_0914_, w_0666_, w_0778_);
not (w_0024_, in10[1]);
or (w_0735_, w_0193_, w_0525_);
and (w_0401_, w_0088_, w_0324_);
not (w_0779_, w_0199_);
and (w_0587_, w_0576_, w_0626_);
not (w_0898_, in10[0]);
or (w_0799_, w_0737_, w_0770_);
or (w_0501_, w_0271_, w_0142_);
and (w_0213_, w_1015_, w_0947_);
or (w_0102_, in1[1], in2[1]);
and (w_0158_, w_0204_, w_0531_);
or (w_0936_, w_0308_, w_0036_);
or (w_0654_, w_0396_, w_0576_);
and (w_0112_, w_0187_, w_0279_);
or (out6[2], w_0337_, w_0742_);
and (w_0082_, w_0980_, w_0132_);
not (w_1013_, w_0668_);
and (w_0360_, w_0193_, w_0525_);
or (w_0798_, w_0820_, w_0760_);
and (w_0865_, w_0662_, w_0263_);
or (w_0953_, in14[2], w_0751_);
or (w_0068_, in11[1], w_0265_);
and (out14[3], w_0577_, w_0225_);
or (w_0854_, w_0517_, w_0049_);
or (w_0569_, w_0353_, w_0126_);
or (w_0139_, in10[3], w_1024_);
and (w_0877_, w_0400_, w_0178_);
and (w_0727_, in14[2], w_0751_);
not (w_0322_, in15[3]);
not (w_0984_, w_0601_);
or (w_0762_, w_0723_, w_0229_);
or (w_0239_, w_0758_, w_0010_);
and (w_0965_, w_0996_, w_1006_);
and (w_0103_, w_0116_, w_0469_);
not (w_0672_, in7[0]);
and (w_0412_, w_0915_, w_0718_);
not (w_0295_, w_0172_);
and (w_0347_, w_1022_, w_0003_);
and (w_0773_, w_0939_, w_0916_);
not (w_0891_, in4[0]);
or (w_0624_, in14[4], w_0262_);
or (w_0237_, w_0930_, w_0565_);
and (w_0542_, w_0970_, w_0802_);
or (w_0869_, w_0719_, w_0965_);
and (w_0719_, w_0148_, w_0958_);
not (w_0317_, in8[1]);
and (w_1015_, w_0915_, w_0901_);
or (w_0003_, w_0397_, w_0837_);
and (w_0978_, w_0835_, w_0354_);
or (w_0195_, w_0058_, w_0065_);
and (w_0337_, w_0033_, w_0534_);
or (w_1011_, w_1003_, w_0327_);
and (w_0979_, w_0554_, w_0974_);
and (w_0929_, w_0986_, w_0647_);
and (w_0638_, w_0388_, w_0414_);
or (w_0766_, w_0015_, w_0052_);
or (w_0514_, w_0164_, w_0357_);
or (w_0459_, w_0561_, w_0387_);
or (w_0795_, w_0945_, w_0958_);
or (w_0382_, w_0989_, w_0659_);
and (w_0753_, w_0323_, w_0707_);
or (w_0738_, w_0727_, w_0127_);
or (w_0093_, w_0120_, w_0782_);
or (w_0995_, w_0011_, w_0482_);
or (w_0284_, w_0897_, w_0711_);
and (w_0463_, w_0210_, w_0664_);
or (w_0521_, w_0381_, w_0827_);
and (w_0677_, w_0073_, w_0043_);
or (w_0186_, w_0854_, w_0344_);
and (w_0688_, in11[1], w_0265_);
or (w_0005_, w_0185_, w_0471_);
or (w_0206_, w_0950_, w_0283_);
or (w_0449_, w_0868_, w_0811_);
or (w_0403_, w_0383_, w_0973_);
and (w_0710_, w_0721_, w_0340_);
not (w_0429_, in6[0]);
or (w_0159_, w_0009_, w_0233_);
and (w_0942_, w_0331_, w_0563_);
or (w_0172_, w_0407_, w_0309_);
not (w_0125_, w_0585_);
or (out13[2], w_0948_, w_0401_);
and (w_0745_, in2[0], w_0280_);
or (w_0171_, w_0331_, w_0563_);
or (w_0985_, w_0836_, w_0282_);
and (w_0920_, w_0989_, w_0924_);
or (w_0575_, w_0236_, w_0222_);
and (w_0661_, w_0641_, w_0911_);
and (w_0123_, w_0775_, w_0488_);
and (w_0204_, w_0776_, w_0464_);
and (w_0489_, w_0755_, w_0644_);
or (w_0700_, w_0588_, w_0276_);
not (w_0517_, in9[0]);
and (out11[0], w_0289_, w_0016_);
or (out7[2], w_0189_, w_0993_);
or (out4[1], w_0201_, w_0971_);
and (w_0616_, w_0765_, w_0683_);
or (w_0191_, w_0773_, w_0252_);
not (w_0106_, w_0630_);
and (w_0090_, in15[1], w_0634_);
or (w_0154_, w_0259_, w_0566_);
and (w_0608_, w_0404_, w_0941_);
or (w_0633_, w_0054_, w_0530_);
or (out5[1], w_0435_, w_0920_);
or (w_0911_, w_0542_, w_0942_);
not (w_0236_, w_0000_);
or (w_0505_, w_0765_, w_0364_);
or (out14[0], w_0722_, w_0105_);
and (w_0561_, w_0118_, w_0569_);
or (w_0718_, w_0512_, w_0673_);
and (w_0440_, in10[1], w_0695_);
or (w_0303_, w_0305_, w_0352_);
and (w_0053_, w_0553_, w_0762_);
or (out12[0], w_0158_, w_0377_);
and (w_0983_, w_0746_, w_0697_);
and (w_0357_, w_0467_, w_0493_);
or (out2[0], w_0572_, w_0788_);
not (w_0367_, w_0840_);
or (w_0858_, w_0712_, w_0103_);
and (w_0684_, w_0215_, w_0508_);
not (w_0937_, w_0068_);
and (w_1001_, w_0420_, w_0819_);
or (w_0909_, w_0020_, w_0548_);
and (w_0653_, w_0402_, w_0862_);
and (w_0160_, w_0878_, w_0617_);
and (w_0895_, w_0270_, w_0652_);
or (w_0903_, in13[3], in12[3]);
or (w_0373_, in10[2], w_0025_);
not (w_0180_, w_0470_);
or (w_0879_, w_0831_, w_0318_);
and (w_0863_, w_0017_, w_0838_);
or (w_0280_, w_0177_, w_0519_);
or (w_0142_, w_0914_, w_0674_);
or (w_0140_, w_0821_, w_0591_);
or (w_0372_, w_0273_, w_0934_);
and (w_0274_, w_0210_, w_0842_);
and (w_0746_, w_0136_, w_0822_);
not (w_0756_, w_0145_);
and (w_0235_, w_0218_, w_0526_);
and (w_0475_, in9[4], in8[4]);
or (w_0736_, w_0402_, w_0862_);
and (w_0361_, w_0083_, w_0121_);
and (w_0371_, in10[0], w_0390_);
and (w_1022_, w_0734_, w_0115_);
or (w_0922_, w_1017_, w_0846_);
or (w_0526_, w_0307_, w_0067_);
not (w_0849_, in8[2]);
or (w_0366_, w_0011_, w_0848_);
and (w_0954_, w_0425_, w_0935_);
and (w_0940_, w_0697_, w_1018_);
and (w_0377_, w_0617_, w_0047_);
not (w_0750_, in14[3]);
or (w_0660_, w_0207_, w_1009_);
not (w_0302_, w_0069_);
or (w_0344_, w_1017_, w_0114_);
or (w_0574_, w_0866_, w_0978_);
and (w_0765_, w_0219_, w_0093_);
and (w_0426_, w_0738_, w_0764_);
not (w_0631_, w_0431_);
or (w_0293_, in14[3], w_0355_);
or (w_0378_, w_0013_, w_0588_);
or (w_0749_, w_0544_, w_0648_);
and (w_0873_, w_0981_, w_0095_);
or (w_0915_, w_0182_, w_0399_);
not (w_0223_, w_0941_);
or (w_0258_, w_0932_, w_0682_);
and (out6[0], w_0080_, w_0527_);
or (w_0692_, w_0079_, w_0700_);
and (w_1017_, in9[1], in8[1]);
not (w_0212_, w_0914_);
and (w_0646_, in13[3], in12[3]);
and (w_0982_, w_0878_, w_0941_);
or (w_0883_, w_0087_, w_0261_);
not (w_0097_, in14[0]);
and (w_0111_, in11[0], w_0061_);
or (w_0479_, w_0869_, w_0642_);
or (w_0531_, w_0647_, w_0987_);
and (w_0230_, w_0171_, w_0094_);
or (w_0441_, w_0017_, w_0838_);
and (w_0273_, in10[2], w_0025_);
or (w_0783_, in6[1], w_0409_);
and (w_0444_, w_0800_, w_0533_);
or (w_0668_, in13[1], in12[1]);
and (w_0427_, w_0592_, w_0583_);
and (w_0545_, w_0294_, w_0847_);
not (w_0062_, in13[1]);
and (w_0405_, w_0259_, w_0566_);
and (w_0175_, w_0363_, w_0803_);
or (out13[0], w_0745_, w_0611_);
not (w_0049_, in8[0]);
or (w_0923_, w_0730_, w_0998_);
and (w_0060_, w_0485_, w_0432_);
or (w_0900_, w_0813_, w_0362_);
or (w_0516_, w_0356_, w_0291_);
and (w_0472_, w_1008_, w_0363_);
and (w_0639_, w_0427_, w_0689_);
and (w_0415_, w_1011_, w_0006_);
or (w_0073_, w_0499_, w_0613_);
or (out1[1], w_0417_, w_0865_);
or (w_0041_, w_0192_, w_0523_);
not (w_0991_, in13[0]);
or (out9[1], w_0109_, w_0619_);
or (w_0663_, w_0716_, w_0128_);
or (w_0439_, in15[2], w_0314_);
and (w_0130_, w_0524_, w_0484_);
not (w_0386_, w_0551_);
and (w_0997_, w_0902_, w_0771_);
or (w_0810_, w_0961_, w_0653_);
and (w_0934_, w_0874_, w_0451_);
or (w_0655_, w_0371_, w_0926_);
and (w_0087_, in15[3], w_0705_);
not (w_0114_, w_0905_);
or (w_0557_, w_0272_, w_0610_);
and (w_1006_, w_0118_, w_0630_);
and (w_0096_, w_0037_, w_0546_);
or (w_0028_, w_0394_, w_0982_);
not (w_0033_, w_0579_);
and (w_0853_, w_0404_, w_0424_);
and (w_1021_, w_0758_, w_0928_);
or (w_0606_, in10[1], w_0695_);
or (w_0219_, w_0104_, w_0476_);
not (w_0499_, in11[4]);
not (w_0375_, w_0903_);
and (w_0835_, w_0413_, w_0458_);
or (w_0838_, w_0482_, w_0448_);
or (w_0395_, w_0220_, w_0816_);
and (w_0418_, w_0972_, w_0736_);
or (out8[2], w_0964_, w_0286_);
or (w_0384_, in13[2], in12[2]);
not (w_0547_, w_0961_);
or (w_0829_, w_0467_, w_0493_);
and (w_0994_, w_0138_, w_0845_);
or (w_1019_, w_0427_, w_0689_);
and (w_1003_, w_0183_, w_0433_);
and (w_0623_, w_0835_, w_1016_);
or (w_0241_, w_0150_, w_0076_);
and (w_0846_, w_0398_, w_0031_);
or (w_0532_, w_0013_, w_0256_);
and (w_0868_, w_0474_, w_0035_);
and (w_0918_, w_1022_, w_0895_);
or (w_0214_, w_0804_, w_0801_);
not (w_0669_, in8[3]);
or (w_0124_, w_0413_, w_0458_);
and (w_0267_, w_0190_, w_0345_);
not (w_0197_, in12[3]);
not (w_0648_, w_0139_);
and (w_0177_, w_0576_, w_0813_);
and (w_0581_, w_0009_, w_0576_);
and (w_0301_, w_0781_, w_0735_);
not (w_0843_, w_0456_);
and (w_0008_, w_0730_, w_0998_);
or (w_0680_, w_0515_, w_0882_);
and (w_0128_, w_0076_, w_0175_);
and (w_0095_, w_0755_, w_0709_);
and (w_0399_, w_0990_, w_0452_);
or (out3[0], w_0999_, w_0063_);
and (w_0430_, w_0472_, w_0879_);
or (w_0333_, w_0220_, w_0412_);
not (w_0776_, w_0977_);
not (w_0777_, w_0443_);
or (w_0541_, w_0514_, w_0765_);
not (w_0266_, w_0390_);
and (w_1018_, w_0864_, w_0506_);
or (w_0925_, w_0411_, w_0912_);
and (w_0878_, w_0856_, w_0628_);
and (w_0352_, w_0528_, w_0167_);
or (w_0893_, w_0608_, w_0785_);
and (w_0682_, w_0244_, w_0288_);
or (w_0679_, in9[0], in8[0]);
and (w_0029_, w_0724_, w_0311_);
and (w_0075_, w_0950_, w_0283_);
or (w_0037_, w_0574_, w_0774_);
or (w_0169_, w_0076_, w_0175_);
or (out11[3], w_0374_, w_0623_);
and (w_0589_, w_0325_, w_0378_);
and (w_0278_, w_0772_, w_0232_);
or (w_0652_, w_0897_, w_0250_);
and (w_0964_, w_0179_, w_0946_);
and (w_0038_, in15[4], w_0808_);
not (w_0921_, w_0739_);
or (w_0803_, w_0502_, w_0066_);
or (w_0793_, w_0491_, w_0328_);
or (w_0591_, w_0727_, w_0078_);
and (w_0643_, w_0980_, w_0209_);
or (w_0247_, in14[0], w_0490_);
and (w_0894_, w_0549_, w_0148_);
or (w_0901_, w_1011_, w_0006_);
or (w_0493_, w_0688_, w_0937_);
and (w_0935_, w_0487_, w_0470_);
and (w_0455_, w_0406_, w_0578_);
or (w_0657_, w_0030_, w_0074_);
or (w_0628_, in3[0], w_0706_);
and (w_1023_, w_0919_, w_0944_);
and (w_0176_, w_0399_, w_0175_);
and (w_0702_, in6[0], w_0892_);
and (w_0764_, w_0423_, w_0293_);
and (w_0085_, w_0945_, w_0129_);
and (w_0805_, w_0148_, w_0758_);
or (w_0339_, w_0593_, w_0010_);
and (w_0436_, w_0917_, w_0627_);
or (w_0772_, w_0351_, w_1020_);
and (w_0926_, w_0543_, w_0606_);
not (w_0051_, w_0124_);
not (w_0645_, w_0265_);
and (w_0861_, w_0967_, w_0237_);
and (w_0354_, w_0793_, w_0349_);
or (w_0107_, in13[0], in12[0]);
or (w_0019_, w_0863_, w_0698_);
or (out9[0], w_0473_, w_0607_);
or (w_0693_, w_0988_, w_0867_);
or (w_0002_, w_0097_, w_0536_);
or (w_0126_, w_0719_, w_0106_);
and (w_0462_, w_0664_, w_0161_);
or (w_0183_, w_0320_, w_0518_);
or (w_0086_, w_0372_, w_0640_);
or (w_0871_, in4[1], in5[1]);
or (w_0358_, w_0039_, w_0123_);
not (w_0058_, w_0244_);
or (w_0508_, in9[2], in8[2]);
and (w_0207_, w_0869_, w_0642_);
and (w_0930_, w_0700_, w_0179_);
and (w_0471_, w_0077_, w_0182_);
or (out13[1], w_0231_, w_0954_);
or (w_0704_, w_0263_, w_0633_);
not (w_0943_, in13[2]);
and (w_0042_, w_0622_, w_0084_);
and (w_0664_, w_0163_, w_0701_);
or (w_0812_, w_0385_, w_0518_);
and (w_0884_, w_0633_, w_0235_);
and (w_0518_, w_0104_, w_0200_);
or (w_0578_, in14[1], w_0230_);
and (w_0141_, w_0237_, w_0697_);
or (w_0094_, w_0970_, w_0802_);
and (w_0325_, w_0064_, w_0443_);
or (w_0423_, w_0750_, w_0693_);
not (w_0715_, w_0904_);
or (out7[1], w_0929_, w_0316_);
or (w_0629_, w_0767_, w_0368_);
and (w_0074_, w_0274_, w_0575_);
not (w_0166_, in11[2]);
or (w_0919_, w_0681_, w_0542_);
not (w_0611_, w_0740_);
or (w_0221_, w_0515_, w_0367_);
or (w_0089_, w_0800_, w_0533_);
and (w_0370_, w_1022_, w_0987_);
or (w_0875_, w_0127_, w_0951_);
or (w_0257_, w_0662_, w_0486_);
and (w_0217_, w_0116_, w_0629_);
or (w_0670_, w_0560_, w_0455_);
or (w_0852_, w_0048_, w_0851_);
not (w_0181_, in13[3]);
or (w_0577_, w_1001_, w_0015_);
or (w_0833_, w_0768_, w_0404_);
or (w_0040_, w_0728_, w_0165_);
not (w_0949_, w_0695_);
and (w_0593_, w_0644_, w_0457_);
and (w_0390_, w_0854_, w_0679_);
and (w_0714_, w_0797_, w_0781_);
not (w_0549_, w_0691_);
and (w_0355_, w_0191_, w_0909_);
and (w_0052_, w_0784_, w_0163_);
and (w_0618_, w_0507_, w_0962_);
or (w_0045_, w_0680_, w_0248_);
and (w_0315_, in3[0], w_0706_);
and (w_0728_, w_0438_, w_0186_);
or (w_0864_, w_0187_, w_0168_);
or (w_0059_, w_0385_, w_0204_);
and (w_0698_, w_0009_, w_0079_);
and (w_0261_, w_0618_, w_0350_);
or (w_0603_, w_0101_, w_0661_);
not (w_0108_, w_0352_);
or (out12[2], w_0587_, w_1021_);
or (w_0709_, w_0774_, w_0746_);
or (w_0904_, in10[4], w_0602_);
and (w_1004_, w_0076_, w_0198_);
and (w_0393_, w_0297_, w_0521_);
and (w_0946_, w_1010_, w_0258_);
and (w_0515_, in11[4], w_0418_);
not (w_0196_, w_0436_);
or (w_0662_, w_0556_, w_0744_);
or (w_0411_, w_0968_, w_0777_);
not (w_0098_, in5[0]);
or (w_0787_, in10[0], w_0390_);
or (w_0443_, in11[3], w_0146_);
and (w_1009_, w_0561_, w_0387_);
and (w_0913_, w_0169_, w_0218_);
or (out5[0], w_0249_, w_1002_);
or (w_0272_, w_0087_, w_0174_);
and (w_0046_, w_0631_, w_0313_);
or (w_0966_, w_0666_, w_0778_);
or (w_0179_, w_0405_, w_0075_);
or (w_0665_, w_0088_, w_0346_);
and (w_0747_, w_0524_, w_0732_);
or (w_0758_, w_0503_, w_0696_);
and (w_0192_, in1[0], in2[0]);
and (w_0599_, w_0385_, w_0204_);
or (w_0967_, w_0586_, w_0612_);
and (w_0199_, w_0257_, w_0570_);
or (w_0962_, in15[3], w_0705_);
or (w_0498_, w_0898_, w_0266_);
and (w_0010_, w_0901_, w_0333_);
not (w_0004_, in4[1]);
and (w_0813_, w_0510_, w_0465_);
and (w_0757_, w_0658_, w_0540_);
and (w_0327_, w_0059_, w_0264_);
and (w_0297_, w_0647_, w_0395_);
and (w_0398_, in9[0], in8[0]);
or (w_0446_, w_0138_, w_0125_);
and (w_0548_, w_0022_, w_0903_);
or (w_0072_, w_0307_, w_0001_);
or (w_0000_, w_0039_, w_0077_);
or (w_0627_, w_0874_, w_0451_);
not (w_0641_, in14[1]);
and (w_0636_, w_0516_, w_0605_);
not (w_0188_, w_0892_);
or (w_0512_, w_0558_, w_0155_);
or (w_0996_, w_0608_, w_0729_);
or (w_0243_, w_0381_, w_0360_);
or (w_0580_, w_0713_, w_0199_);
and (out11[2], w_0026_, w_0960_);
or (w_0200_, in7[0], w_0994_);
not (w_0806_, w_0200_);
and (w_0253_, w_0307_, w_0067_);
and (w_0353_, w_0194_, w_0487_);
and (w_0174_, w_0322_, w_0131_);
or (w_0842_, w_0784_, w_0485_);
and (w_0523_, w_0756_, w_0102_);
not (w_0848_, w_0044_);
or (w_0167_, in9[3], in8[3]);
and (w_0573_, w_0700_, w_0021_);
and (w_0808_, w_0214_, w_0089_);
not (w_0790_, in12[2]);
or (w_0209_, w_0776_, w_0152_);
not (w_0296_, w_0706_);
and (w_0318_, w_0028_, w_0123_);
and (w_0157_, w_0353_, w_0126_);
or (w_0950_, w_0639_, w_0278_);
or (w_0104_, w_0672_, w_0731_);
not (w_0613_, w_0418_);
and (w_0047_, w_0453_, w_0251_);
not (w_0520_, in5[1]);
or (w_0092_, w_0360_, w_0393_);
not (w_0468_, w_0373_);
or (w_0786_, w_0922_, w_0684_);
and (w_0466_, w_0804_, w_0801_);
and (w_0963_, w_0182_, w_0399_);
and (w_0265_, w_0478_, w_0655_);
or (w_0012_, w_0222_, w_0361_);
or (w_0026_, w_0601_, w_0419_);
or (w_0244_, w_0148_, w_0987_);
and (w_0582_, in6[1], w_0409_);
and (w_0656_, w_0560_, w_0455_);
or (w_0972_, w_0877_, w_0149_);
and (w_0077_, w_0654_, w_0202_);
or (w_0845_, in6[0], w_0892_);
and (w_0381_, w_0593_, w_0010_);
or (w_0730_, w_0038_, w_0832_);
or (w_0227_, in4[0], in5[0]);
or (out14[1], w_0275_, w_0463_);
or (w_0270_, w_0323_, w_0005_);
or (w_0701_, w_0407_, w_0147_);
or (w_0712_, w_0185_, w_0959_);
not (w_0761_, in12[1]);
and (w_0442_, w_0574_, w_0774_);
or (w_0203_, w_0772_, w_0232_);
and (w_0242_, w_0017_, w_0758_);
or (w_0084_, w_0537_, w_0815_);
and (w_0816_, w_1003_, w_0327_);
or (w_0957_, w_0273_, w_0468_);
or (w_0952_, w_0700_, w_0179_);
or (w_0769_, w_0919_, w_0944_);
or (w_0691_, w_0914_, w_0008_);
and (w_0055_, w_0712_, w_0103_);
and (w_0263_, w_0829_, w_0889_);
and (w_0310_, w_0774_, w_0746_);
and (w_1014_, w_0220_, w_0412_);
or (w_0163_, w_0039_, w_0489_);
and (w_0481_, w_0714_, w_0226_);
and (w_0145_, in1[1], in2[1]);
and (w_0032_, w_0224_, w_0240_);
and (w_0782_, w_0382_, w_0596_);
or (w_0264_, w_0878_, w_0617_);
and (w_0844_, w_0022_, w_0191_);
and (w_0069_, w_0592_, w_0871_);
or (w_0820_, w_0968_, w_0589_);
and (w_0821_, w_0406_, w_0686_);
or (w_0034_, w_0454_, w_0927_);
or (w_0778_, w_0571_, w_0444_);
not (w_0989_, in7[1]);
or (w_0433_, w_0224_, w_0524_);
or (w_0406_, w_0641_, w_0911_);
or (w_0043_, w_0796_, w_0221_);
and (w_0283_, w_0382_, w_0219_);
or (w_0368_, w_0861_, w_0060_);
or (w_1008_, w_0432_, w_1022_);
or (w_0289_, w_0385_, w_0083_);
and (w_0910_, w_0034_, w_0175_);
and (w_0742_, w_0579_, w_0888_);
and (w_0013_, in11[2], w_0436_);
and (w_0823_, w_0091_, w_0504_);
or (w_0724_, w_0141_, w_0359_);
and (w_0245_, in1[1], w_0173_);
and (w_0153_, w_0767_, w_0368_);
or (w_0504_, in11[2], w_0436_);
and (w_0759_, w_0977_, w_0082_);
and (w_0348_, w_0878_, w_0524_);
and (w_0737_, w_0037_, w_0057_);
and (w_0706_, w_0665_, w_0509_);
or (w_0658_, w_0034_, w_0175_);
and (w_0304_, w_0002_, w_0603_);
or (out4[0], w_0649_, w_0130_);
or (w_0630_, w_0148_, w_0958_);
or (w_0859_, in11[0], w_0061_);
or (w_0938_, w_0440_, w_0635_);
and (w_0291_, w_0305_, w_0352_);
or (w_0134_, w_0474_, w_0035_);
or (w_0870_, w_0062_, w_0761_);
or (w_0734_, w_0009_, w_0576_);
and (w_0987_, w_0376_, w_0890_);
and (w_0642_, w_0843_, w_0814_);
and (w_0927_, w_0039_, w_0489_);
and (w_0959_, w_0897_, w_0250_);
and (w_0397_, w_0050_, w_0956_);
and (w_0559_, w_0237_, w_0673_);
not (w_0822_, w_0982_);
or (out12[1], w_0422_, w_0741_);
and (w_0105_, w_0172_, w_0593_);
and (w_0530_, w_0104_, w_0476_);
or (w_0720_, w_0784_, w_0163_);
or (w_0438_, w_0604_, w_0317_);
and (w_0454_, w_0407_, w_0147_);
or (w_0193_, w_0453_, w_0597_);
or (w_0464_, in15[0], w_0824_);
and (w_0435_, in7[1], w_0370_);
and (w_0342_, w_0192_, w_0523_);
not (w_0632_, w_0409_);
or (w_0168_, w_0708_, w_0392_);
and (w_0687_, in13[4], in12[4]);
or (w_0814_, w_0079_, w_0768_);
or (w_0792_, w_0554_, w_0876_);
or (w_0992_, w_1005_, w_0108_);
and (w_0832_, w_0883_, w_0437_);
or (w_0285_, w_0404_, w_0161_);
or (w_0149_, w_0961_, w_0715_);
and (w_0948_, in1[0], w_0335_);
and (w_0081_, w_0697_, w_0763_);
not (w_0391_, w_0025_);
and (w_0760_, w_0073_, w_0840_);
or (w_0020_, w_0537_, w_1023_);
and (w_1002_, w_0672_, w_0389_);
and (w_0379_, in14[3], w_0355_);
not (w_0137_, in11[3]);
and (w_0259_, w_0203_, w_1019_);
and (w_0999_, w_0434_, w_0284_);
and (w_0182_, w_0541_, w_0704_);
or (w_0840_, in11[4], w_0418_);
and (w_0324_, w_0569_, w_0538_);
not (w_0488_, w_1004_);
and (w_0122_, w_0535_, w_0766_);
or (w_0215_, w_0726_, w_0849_);
and (w_0432_, w_0900_, w_0952_);
and (w_0437_, w_0365_, w_0850_);
or (w_0539_, w_0621_, w_0069_);
and (w_0450_, w_0271_, w_0142_);
and (out6[1], w_0841_, w_0494_);
or (w_0254_, w_0576_, w_0434_);
or (w_0780_, w_0050_, w_0880_);
or (w_0281_, w_0074_, w_0144_);
or (out14[2], w_0122_, w_0096_);
or (w_0980_, w_0294_, w_0847_);
or (w_0857_, w_0688_, w_0164_);
or (w_0596_, in7[1], w_0860_);
and (w_0899_, w_0528_, w_0992_);
not (w_0754_, w_0958_);
not (w_0667_, in10[3]);
and (w_0120_, in7[0], w_0994_);
and (w_0881_, w_0320_, w_0518_);
or (w_0305_, w_0246_, w_0513_);
or (w_0775_, w_0076_, w_0198_);
or (w_0673_, w_0085_, w_0975_);
and (w_0482_, w_0680_, w_0248_);
and (w_0571_, in14[4], w_0262_);
and (w_0079_, w_0349_, w_0045_);
or (w_0707_, w_0986_, w_0554_);
not (w_0408_, w_0298_);
not (w_0651_, in6[1]);
and (w_0109_, w_0945_, w_0205_);
or (w_0452_, w_0945_, w_0129_);
and (w_0428_, w_0750_, w_0693_);
or (w_0396_, w_0832_, w_0598_);
and (out11[1], w_0826_, w_0580_);
or (w_0836_, w_0101_, w_0656_);
and (w_0584_, w_0480_, w_0917_);
and (w_0968_, in11[3], w_0146_);
or (out8[1], w_0616_, w_0884_);
and (w_0537_, in13[2], in12[2]);
not (w_0785_, w_0334_);
and (w_0416_, in7[1], w_0860_);
or (w_0797_, w_0338_, w_0434_);
and (w_0609_, w_0407_, w_0986_);
not (w_0807_, in10[2]);
and (w_0410_, w_0175_, w_0895_);
or (w_0486_, w_0260_, w_0030_);
and (w_0121_, w_0650_, w_0376_);
not (w_0113_, w_0605_);
or (w_0298_, w_0977_, w_0082_);
and (w_0560_, in14[0], w_0490_);
and (w_0851_, w_0969_, w_0439_);
or (w_0647_, w_0055_, w_0153_);
or (w_0889_, w_0111_, w_0341_);
or (w_0685_, w_0444_, w_0466_);
or (w_0022_, w_0181_, w_0197_);
and (w_0827_, w_0338_, w_0434_);
or (w_0323_, w_0123_, w_1003_);
and (w_0619_, w_0662_, w_0983_);
and (w_0224_, w_0467_, w_0859_);
or (w_0527_, w_0224_, w_0941_);
not (w_0495_, in12[0]);
or (w_0309_, w_0805_, w_0896_);
or (w_0990_, w_0662_, w_0198_);
or (w_0876_, w_0160_, w_0599_);
and (w_0017_, w_0690_, w_0124_);
not (w_0815_, w_0384_);
or (w_0590_, w_0398_, w_0031_);
and (w_0598_, w_0676_, w_0023_);
not (w_0511_, in1[1]);
or (w_0818_, w_0729_, w_0180_);
or (w_0292_, w_0516_, w_0605_);
and (w_0741_, w_0129_, w_0703_);
or (w_0385_, w_0315_, w_0564_);
or (w_0683_, w_0253_, w_0595_);
not (w_0690_, w_0835_);
and (w_0722_, w_0295_, w_0338_);
and (w_0232_, w_0326_, w_0446_);
or (w_0334_, w_0404_, w_0941_);
and (w_0231_, in2[1], w_0818_);
or (w_0494_, w_0156_, w_0710_);
and (w_0362_, w_0206_, w_0154_);
and (w_0699_, w_0997_, w_0028_);
not (w_0425_, in2[1]);
and (w_0282_, w_0936_, w_0953_);
or (w_0414_, w_0379_, w_0428_);
or (w_0233_, w_0535_, w_0442_);
and (w_0351_, in4[1], in5[1]);
and (w_0912_, w_0091_, w_0510_);
and (w_0958_, w_0043_, w_0798_);
and (w_0550_, w_0555_, w_0829_);
and (w_0431_, in3[1], w_0071_);
not (w_0099_, w_0464_);
or (w_0136_, w_0878_, w_0941_);
and (w_0148_, w_0885_, w_0594_);
or (w_1010_, w_0913_, w_0195_);
or (w_0152_, w_0090_, w_0545_);
and (w_0497_, in15[2], w_0314_);
and (w_0751_, w_0916_, w_0769_);
and (w_0015_, w_0019_, w_0454_);
or (w_0480_, w_0807_, w_0391_);
and (w_0558_, w_0263_, w_0633_);
and (w_0860_, w_0446_, w_0725_);
not (w_0328_, w_0810_);
and (w_0974_, w_0812_, w_0290_);
not (w_0625_, w_0342_);
and (w_0162_, w_0263_, w_0092_);
or (w_0400_, w_0667_, w_1000_);
and (w_0332_, w_0018_, w_0875_);
or (w_0268_, w_0077_, w_0182_);
or (out13[3], w_0245_, w_0855_);
not (w_0419_, w_0184_);
and (w_0568_, w_1003_, w_0886_);
and (w_0988_, w_0020_, w_0548_);
or (w_0467_, w_0336_, w_0110_);
and (w_0732_, w_0239_, w_0254_);
or (w_0350_, w_0497_, w_0503_);
and (w_0246_, in9[2], in8[2]);
and (w_0066_, w_1008_, w_0117_);
not (w_0771_, w_0894_);
and (w_0788_, w_0399_, w_0112_);
or (w_0313_, in3[1], w_0071_);
or (w_0678_, w_0838_, w_0813_);
or (w_0540_, w_0664_, w_0161_);
not (w_0809_, w_0556_);
and (w_0321_, w_0079_, w_0700_);
or (w_0650_, w_0028_, w_0123_);
not (w_0733_, w_0775_);
and (w_0071_, w_0625_, w_0041_);
not (w_0118_, w_0719_);
or (w_0492_, w_0758_, w_0700_);
or (w_0476_, w_0416_, w_0014_);
and (w_0804_, w_0423_, w_0329_);
and (w_0054_, w_0120_, w_0782_);
and (w_0676_, w_0507_, w_0557_);
and (w_0228_, w_0194_, w_0334_);
and (w_0307_, w_0576_, w_0434_);
and (w_0866_, w_0690_, w_0995_);
and (w_0828_, w_0512_, w_0673_);
or (w_0960_, w_0984_, w_0184_);
and (w_0708_, w_0813_, w_0129_);
and (w_0255_, w_0543_, w_0478_);
or (w_0721_, w_0754_, w_0514_);
not (w_0825_, in3[0]);
or (w_0752_, w_0432_, w_0129_);
or (w_0538_, w_0996_, w_1006_);
or (w_0076_, w_0261_, w_0386_);
and (w_0184_, w_0159_, w_0933_);
or (w_0070_, w_0315_, w_0046_);
and (w_0610_, w_0969_, w_0460_);
or (w_0129_, w_0759_, w_0408_);
and (w_0998_, w_0212_, w_0966_);
or (out9[2], w_0872_, w_1007_);
not (w_0931_, w_0814_);
or (w_0445_, w_0497_, w_0332_);
and (w_0001_, w_0758_, w_0010_);
or (w_0939_, w_0943_, w_0790_);
or (w_0874_, w_0440_, w_0119_);
and (w_0127_, w_0836_, w_0282_);
or (w_0483_, w_0687_, w_0921_);
and (w_0811_, w_0844_, w_0483_);
not (w_0971_, w_0505_);
or (w_0007_, w_0813_, w_0129_);
or (w_0474_, w_0646_, w_0988_);
and (w_0586_, w_0150_, w_0076_);
or (w_0801_, w_0571_, w_0600_);
and (w_0897_, w_0986_, w_0554_);
or (w_0290_, w_0878_, w_0524_);
and (w_0824_, w_0002_, w_0247_);
and (w_0892_, w_0694_, w_0227_);
or (w_0885_, w_0676_, w_0023_);
or (w_0856_, w_0825_, w_0296_);
or (w_0116_, w_0485_, w_0432_);
and (w_0830_, w_0243_, w_0757_);
or (w_0161_, w_0359_, w_0213_);
not (w_0908_, in15[4]);
or (w_0689_, w_0582_, w_0211_);
or (w_0252_, w_0646_, w_0375_);
not (w_0374_, w_0135_);
or (w_0210_, w_0019_, w_0967_);
and (w_0711_, w_0123_, w_1003_);
or (w_0583_, w_0694_, w_0302_);
or (w_0080_, w_0320_, w_0223_);
and (w_0880_, w_0514_, w_0617_);
and (w_0025_, w_0040_, w_0786_);
or (out12[3], w_0853_, w_0208_);
and (w_0485_, w_0833_, w_0241_);
or (w_0551_, w_0618_, w_0350_);
and (w_0867_, w_0773_, w_0252_);
and (w_0061_, w_0498_, w_0787_);
or (w_0594_, w_0883_, w_0437_);
and (w_0579_, w_0721_, w_0841_);
or (out2[1], w_0940_, w_0347_);
or (w_0364_, w_0758_, w_0028_);
and (w_0605_, w_0369_, w_0615_);
or (w_0402_, w_0544_, w_0834_);
not (w_0731_, w_0994_);
or (w_0528_, w_0500_, w_0669_);
or (w_0251_, w_0029_, w_0430_);
and (w_0031_, w_0438_, w_0905_);
or (w_0365_, w_0908_, w_0685_);
or (w_0543_, w_0024_, w_0949_);
or (w_0675_, w_0297_, w_0100_);
and (w_0100_, w_0453_, w_0597_);
and (w_0448_, w_0677_, w_0366_);
and (w_0944_, w_0939_, w_0384_);
or (w_0178_, w_0584_, w_0749_);
and (w_0622_, w_0870_, w_0171_);
and (w_0614_, w_0514_, w_0301_);
or (w_0117_, w_0237_, w_0697_);
not (w_0907_, w_0143_);
and (w_0249_, in7[0], w_0176_);
or (w_0225_, w_0574_, w_0720_);
or (w_0487_, w_0492_, w_0893_);
and (w_0220_, w_0554_, w_0876_);
not (w_0491_, w_0477_);
or (w_0115_, w_0017_, w_0758_);
and (w_0453_, w_0629_, w_0858_);
or (w_0496_, w_0019_, w_0454_);
and (w_0882_, w_0820_, w_0760_);
not (w_0404_, w_0076_);
and (w_0597_, w_1011_, w_0792_);
or (w_0016_, w_0878_, w_0723_);
or (w_0009_, w_0835_, w_0051_);
or (w_0592_, w_0004_, w_0520_);
or (w_0902_, w_0549_, w_0148_);
not (w_0133_, w_0902_);
or (out7[0], w_0081_, w_0918_);
or (w_0886_, w_0348_, w_0839_);
or (w_0319_, w_0309_, w_0512_);
or (w_0387_, w_0456_, w_0931_);
and (w_0621_, in4[0], in5[0]);
and (w_0189_, w_0309_, w_0338_);
or (w_0326_, w_0651_, w_0632_);
not (w_0696_, w_0852_);
not (w_0635_, w_0606_);
not (w_0014_, w_0596_);
or (w_0524_, w_0120_, w_0806_);
and (w_0770_, w_0842_, w_0190_);
and (w_0417_, w_0945_, w_0514_);
not (w_0789_, w_0146_);
and (w_0612_, w_0768_, w_0404_);
and (w_0649_, w_0518_, w_0752_);
endmodule

module sub_module3(
    input wire [2:0] in1,
    input wire [2:0] in2,
    input wire [2:0] in3,
    input wire [3:0] in4,
    input wire [3:0] in5,
    input wire [3:0] in6,
    input wire [4:0] in7,
    input wire [4:0] in8,
    input wire [4:0] in9,
    input wire [5:0] in10,
    input wire [5:0] in11,
    input wire [5:0] in12,
    input wire [6:0] in13,
    input wire [6:0] in14,
    input wire [6:0] in15,
    output wire [1:0] out1,
    output wire [1:0] out2,
    output wire [1:0] out3,
    output wire [1:0] out4,
    output wire [1:0] out5,
    output wire [1:0] out6,
    output wire [1:0] out7,
    output wire [1:0] out8,
    output wire [2:0] out9,
    output wire [2:0] out10,
    output wire [2:0] out11,
    output wire [2:0] out12,
    output wire [2:0] out13,
    output wire [2:0] out14
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
wire w_0945_;
wire w_0946_;
wire w_0947_;
wire w_0948_;
wire w_0949_;
wire w_0950_;
and (w_0403_, w_0727_, w_0486_);
and (w_0187_, w_0727_, w_0083_);
or (w_0775_, in9[3], w_0698_);
and (w_0444_, w_0189_, w_0328_);
or (w_0719_, w_0457_, w_0944_);
or (w_0408_, w_0007_, w_0398_);
or (w_0574_, w_0799_, w_0113_);
or (w_0454_, w_0909_, w_0082_);
or (w_0394_, in9[4], w_0943_);
or (w_0323_, w_0868_, w_0318_);
or (w_0312_, w_0077_, w_0927_);
and (w_0824_, w_0145_, w_0181_);
or (w_0813_, w_0286_, w_0247_);
not (w_0892_, in10[0]);
or (w_0109_, w_0022_, w_0320_);
or (w_0784_, w_0438_, w_0887_);
and (w_0869_, in4[1], in5[1]);
not (w_0269_, in6[1]);
or (w_0003_, w_0727_, w_0486_);
or (w_0537_, w_0836_, w_0048_);
and (out9[0], w_0376_, w_0404_);
or (w_0061_, in4[0], in5[0]);
or (w_0758_, w_0384_, w_0738_);
or (w_0052_, w_0668_, w_0157_);
not (w_0411_, w_0741_);
or (w_0265_, w_0876_, w_0185_);
not (w_0700_, w_0083_);
not (w_0330_, w_0774_);
or (w_0374_, w_0675_, w_0688_);
or (w_0174_, in4[3], in5[3]);
and (w_0034_, w_0261_, w_0409_);
or (w_0250_, w_0658_, w_0463_);
or (w_0786_, w_0261_, w_0043_);
not (w_0932_, in15[1]);
not (w_0388_, in11[2]);
or (w_0793_, w_0089_, w_0900_);
or (w_0768_, w_0247_, w_0096_);
or (out14[0], w_0825_, w_0370_);
or (w_0119_, w_0172_, w_0466_);
and (w_0400_, w_0412_, w_0085_);
and (w_0208_, w_0111_, w_0669_);
and (w_0725_, w_0747_, w_0546_);
and (w_0941_, in12[2], w_0391_);
or (w_0595_, w_0376_, w_0841_);
or (w_0919_, in7[1], in8[1]);
and (w_0621_, w_0330_, w_0743_);
not (w_0135_, in15[2]);
or (w_0045_, w_0086_, w_0874_);
not (w_0228_, w_0506_);
or (w_0555_, in10[3], in11[3]);
and (w_0325_, w_0624_, w_0377_);
and (w_0649_, w_0818_, w_0453_);
and (w_0800_, w_0635_, w_0079_);
not (w_0715_, w_0796_);
not (w_0470_, w_0001_);
and (w_0458_, w_0732_, w_0503_);
or (w_0272_, w_0717_, w_0433_);
not (w_0740_, w_0129_);
or (w_0220_, w_0920_, w_0860_);
or (w_0622_, w_0214_, w_0331_);
and (w_0791_, w_0367_, w_0862_);
and (w_0896_, w_0808_, w_0327_);
and (w_0809_, w_0471_, w_0458_);
or (w_0583_, w_0261_, w_0049_);
and (w_0426_, w_0659_, w_0687_);
or (w_0546_, out4[0], w_0930_);
or (w_0355_, w_0032_, w_0258_);
or (w_0853_, w_0292_, w_0055_);
and (w_0856_, w_0861_, w_0191_);
and (w_0410_, in7[4], in8[4]);
and (w_0098_, w_0660_, w_0859_);
not (w_0048_, in8[1]);
and (w_0874_, w_0607_, w_0721_);
and (w_0590_, w_0541_, w_0821_);
not (w_0877_, w_0935_);
and (w_0744_, w_0842_, w_0858_);
or (w_0138_, in15[5], w_0519_);
or (w_0521_, w_0237_, w_0016_);
and (w_0010_, w_0938_, w_0408_);
and (w_0599_, w_0547_, w_0127_);
or (w_0806_, w_0251_, w_0316_);
or (w_0302_, w_0441_, w_0885_);
or (w_0773_, w_0864_, w_0058_);
and (w_0224_, in13[3], in14[3]);
or (w_0832_, w_0523_, w_0359_);
or (w_0455_, w_0786_, w_0653_);
and (w_0530_, w_0866_, w_0657_);
and (w_0058_, w_0718_, w_0935_);
and (w_0106_, w_0387_, w_0358_);
and (w_0587_, w_0294_, w_0785_);
or (w_0071_, w_0187_, w_0680_);
and (w_0849_, in13[5], in14[5]);
or (w_0328_, w_0611_, w_0312_);
not (w_0532_, w_0896_);
not (w_0385_, w_0003_);
or (w_0209_, w_0634_, w_0341_);
and (w_0847_, w_0793_, w_0589_);
and (w_0831_, w_0406_, w_0649_);
not (w_0210_, w_0687_);
and (w_0675_, in13[2], in14[2]);
or (w_0303_, w_0307_, w_0459_);
or (w_0298_, w_0548_, w_0235_);
or (w_0624_, w_0187_, w_0436_);
or (w_0069_, w_0231_, w_0812_);
and (w_0873_, w_0583_, w_0149_);
or (w_0294_, w_0710_, w_0429_);
and (w_0151_, w_0095_, w_0845_);
and (w_0654_, w_0835_, w_0065_);
or (out10[0], w_0321_, w_0282_);
or (w_0488_, w_0631_, w_0615_);
or (w_0925_, w_0276_, w_0091_);
and (w_0129_, w_0612_, w_0128_);
and (w_0457_, w_0776_, w_0735_);
or (w_0835_, w_0295_, w_0798_);
or (w_0222_, w_0913_, w_0344_);
or (out8[1], w_0863_, w_0297_);
and (w_0860_, in9[3], w_0698_);
or (w_0318_, w_0940_, w_0809_);
and (w_0124_, w_0539_, w_0046_);
and (w_0846_, w_0417_, w_0555_);
not (w_0891_, in14[3]);
not (w_0389_, w_0261_);
or (w_0201_, w_0357_, w_0036_);
or (w_0300_, w_0508_, w_0402_);
or (w_0499_, w_0218_, w_0663_);
not (w_0564_, in14[5]);
not (w_0895_, w_0439_);
and (w_0285_, w_0332_, w_0763_);
and (w_0273_, w_0362_, w_0192_);
not (w_0217_, w_0758_);
not (w_0397_, in5[0]);
and (w_0519_, w_0638_, w_0906_);
and (w_0256_, w_0757_, w_0606_);
not (w_0334_, w_0034_);
or (w_0562_, w_0288_, w_0796_);
and (w_0648_, w_0806_, w_0363_);
not (w_0152_, in5[1]);
or (w_0313_, w_0618_, w_0746_);
and (w_0038_, w_0913_, w_0240_);
not (w_0468_, w_0171_);
not (w_0356_, in4[0]);
or (w_0475_, w_0629_, w_0035_);
or (w_0794_, w_0861_, w_0191_);
or (w_0854_, w_0406_, w_0761_);
or (out6[1], w_0090_, w_0518_);
and (w_0202_, w_0060_, w_0921_);
and (w_0412_, w_0679_, w_0476_);
or (w_0529_, w_0693_, w_0273_);
not (w_0245_, w_0192_);
and (w_0883_, w_0679_, w_0725_);
or (w_0105_, w_0762_, w_0643_);
and (w_0117_, w_0931_, w_0317_);
or (w_0198_, w_0666_, w_0592_);
or (w_0662_, w_0145_, w_0181_);
and (w_0043_, w_0548_, w_0235_);
and (w_0428_, w_0607_, w_0239_);
or (w_0483_, w_0931_, w_0317_);
and (w_0251_, in7[1], in8[1]);
and (w_0482_, w_0159_, w_0880_);
and (w_0825_, w_0755_, w_0431_);
and (w_0902_, w_0775_, w_0828_);
and (w_0023_, w_0570_, w_0175_);
and (w_0057_, w_0322_, w_0024_);
and (w_0661_, in9[2], w_0226_);
and (w_0943_, w_0934_, w_0383_);
and (w_0268_, w_0727_, w_0193_);
and (w_0717_, in12[4], w_0830_);
and (w_0364_, in3[1], w_0464_);
and (w_0685_, w_0073_, w_0150_);
or (w_0168_, w_0206_, w_0026_);
and (w_0884_, w_0417_, w_0612_);
or (w_0552_, w_0849_, w_0496_);
or (w_0718_, w_0437_, w_0098_);
and (w_0930_, w_0497_, w_0644_);
or (w_0088_, w_0480_, w_0618_);
not (w_0802_, in12[1]);
or (w_0176_, w_0499_, w_0850_);
or (w_0219_, w_0908_, w_0857_);
not (w_0513_, w_0308_);
not (w_0502_, w_0464_);
and (w_0745_, w_0241_, w_0380_);
not (w_0159_, w_0130_);
and (w_0422_, w_0235_, w_0504_);
and (w_0270_, w_0374_, w_0027_);
or (w_0876_, w_0939_, w_0534_);
and (out2[0], w_0201_, w_0165_);
not (w_0314_, w_0410_);
or (w_0104_, w_0356_, w_0397_);
and (w_0565_, w_0835_, w_0818_);
or (w_0731_, w_0727_, w_0193_);
not (w_0637_, in13[4]);
or (w_0099_, w_0879_, w_0867_);
and (w_0505_, w_0750_, w_0199_);
or (w_0821_, in10[0], in11[0]);
or (w_0783_, w_0062_, w_0280_);
or (w_0304_, w_0197_, w_0281_);
or (w_0192_, in1[1], in2[1]);
or (w_0931_, w_0325_, w_0435_);
or (w_0083_, w_0422_, w_0873_);
not (w_0145_, w_0351_);
and (out4[1], w_0686_, w_0913_);
or (w_0036_, w_0826_, w_0339_);
not (w_0501_, w_0384_);
or (w_0366_, w_0889_, w_0895_);
not (w_0213_, in4[2]);
not (w_0528_, w_0812_);
or (w_0423_, w_0446_, w_0527_);
and (w_0301_, w_0911_, w_0765_);
not (w_0243_, w_0843_);
not (w_0948_, w_0146_);
not (w_0776_, w_0187_);
not (w_0491_, w_0257_);
and (w_0605_, w_0357_, w_0914_);
and (w_0548_, w_0773_, w_0396_);
or (out13[2], w_0500_, w_0215_);
or (w_0167_, w_0568_, w_0701_);
or (w_0950_, w_0678_, w_0092_);
and (w_0728_, w_0868_, w_0318_);
or (w_0636_, w_0480_, w_0249_);
not (w_0647_, w_0018_);
and (w_0940_, w_0355_, w_0820_);
or (w_0938_, w_0541_, w_0029_);
or (w_0040_, w_0725_, w_0313_);
or (out3[0], w_0759_, w_0023_);
or (w_0238_, w_0823_, w_0124_);
or (w_0866_, w_0444_, w_0730_);
or (w_0545_, w_0526_, w_0751_);
not (w_0751_, w_0079_);
or (w_0601_, w_0285_, w_0283_);
or (w_0730_, w_0509_, w_0025_);
not (w_0707_, in11[0]);
not (w_0420_, w_0396_);
or (w_0332_, w_0274_, w_0032_);
or (w_0689_, w_0838_, w_0564_);
and (w_0320_, w_0301_, w_0205_);
not (w_0399_, w_0864_);
or (w_0487_, w_0263_, w_0915_);
not (out1[0], w_0570_);
and (w_0307_, w_0353_, w_0949_);
not (w_0912_, w_0733_);
or (w_0126_, w_0364_, w_0520_);
and (w_0193_, w_0450_, w_0094_);
and (w_0608_, w_0619_, w_0673_);
and (w_0680_, w_0562_, w_0700_);
or (w_0311_, w_0941_, w_0255_);
not (w_0769_, w_0268_);
or (w_0441_, w_0717_, w_0144_);
and (w_0609_, w_0018_, w_0488_);
and (w_0879_, w_0911_, w_0692_);
not (w_0705_, in1[0]);
and (w_0378_, w_0776_, w_0947_);
and (w_0631_, w_0679_, w_0254_);
and (w_0535_, in12[5], w_0608_);
and (w_0826_, in6[0], w_0817_);
and (w_0016_, w_0153_, w_0136_);
and (w_0908_, in12[3], w_0129_);
or (w_0597_, w_0659_, w_0816_);
or (w_0671_, w_0100_, w_0896_);
or (w_0672_, w_0628_, w_0585_);
not (w_0204_, w_0267_);
not (w_0900_, w_0830_);
and (w_0437_, in4[2], in5[2]);
and (w_0372_, w_0672_, w_0053_);
and (w_0235_, w_0389_, w_0950_);
or (w_0465_, in7[2], in8[2]);
and (w_0827_, w_0689_, w_0308_);
not (w_0435_, w_0580_);
and (w_0349_, w_0351_, w_0229_);
and (w_0137_, w_0791_, w_0207_);
or (w_0194_, w_0642_, w_0714_);
or (w_0143_, w_0530_, w_0579_);
and (w_0321_, w_0583_, w_0050_);
or (w_0184_, w_0279_, w_0601_);
and (w_0496_, w_0489_, w_0827_);
and (w_0588_, w_0791_, w_0303_);
or (w_0490_, w_0565_, w_0340_);
and (w_0646_, w_0712_, w_0116_);
not (w_0682_, w_0280_);
and (w_0170_, w_0214_, w_0331_);
not (w_0240_, w_0473_);
not (w_0218_, w_0876_);
and (w_0466_, w_0442_, w_0002_);
or (w_0694_, w_0354_, w_0336_);
and (w_0258_, w_0183_, w_0494_);
or (w_0571_, w_0913_, w_0240_);
or (w_0262_, w_0216_, w_0006_);
not (w_0814_, w_0072_);
or (w_0424_, w_0617_, w_0118_);
or (w_0514_, w_0478_, w_0223_);
or (w_0497_, w_0607_, w_0721_);
or (w_0232_, w_0084_, w_0097_);
and (w_0709_, w_0584_, w_0543_);
or (w_0072_, w_0605_, w_0291_);
not (w_0651_, w_0043_);
not (w_0339_, w_0563_);
and (w_0230_, in13[4], in14[4]);
and (w_0737_, w_0406_, w_0761_);
or (w_0906_, w_0489_, w_0827_);
and (w_0567_, w_0854_, w_0602_);
and (w_0526_, w_0362_, w_0787_);
and (out13[1], w_0076_, w_0304_);
and (w_0805_, w_0294_, w_0163_);
or (w_0547_, w_0239_, w_0530_);
not (w_0134_, in2[1]);
and (w_0223_, w_0497_, w_0747_);
or (w_0028_, w_0520_, w_0805_);
not (w_0591_, in15[3]);
and (w_0542_, w_0177_, w_0899_);
or (w_0947_, w_0727_, w_0083_);
or (w_0569_, w_0286_, w_0903_);
or (w_0687_, in15[0], w_0115_);
and (w_0347_, w_0790_, w_0945_);
or (w_0898_, in15[3], w_0729_);
or (out9[2], w_0482_, w_0594_);
not (w_0581_, w_0136_);
or (w_0053_, w_0073_, w_0150_);
and (w_0553_, w_0313_, w_0030_);
and (w_0085_, w_0602_, w_0323_);
not (w_0271_, w_0315_);
and (w_0081_, w_0772_, w_0365_);
and (w_0286_, in13[6], in14[6]);
or (w_0365_, w_0629_, w_0470_);
or (w_0246_, w_0894_, w_0481_);
not (w_0075_, w_0116_);
and (w_0015_, in7[3], in8[3]);
or (w_0478_, w_0588_, w_0186_);
and (w_0743_, w_0468_, w_0146_);
not (w_0795_, in13[3]);
or (w_0367_, w_0290_, w_0311_);
or (w_0764_, w_0338_, w_0646_);
or (w_0677_, in1[2], in2[2]);
or (w_0580_, w_0624_, w_0377_);
and (w_0352_, w_0222_, w_0040_);
or (w_0669_, w_0254_, w_0083_);
or (w_0695_, w_0294_, w_0163_);
or (w_0253_, w_0902_, w_0220_);
or (w_0146_, w_0199_, w_0473_);
not (w_0863_, w_0143_);
or (w_0558_, w_0031_, w_0013_);
or (w_0946_, w_0344_, w_0028_);
not (w_0173_, w_0483_);
and (w_0382_, w_0176_, w_0204_);
and (w_0310_, w_0767_, w_0105_);
and (w_0686_, w_0194_, w_0764_);
or (w_0315_, in6[2], w_0361_);
not (w_0568_, w_0376_);
not (w_0890_, w_0773_);
or (w_0471_, w_0588_, w_0288_);
or (w_0131_, w_0758_, w_0368_);
and (w_0123_, w_0837_, w_0652_);
or (w_0158_, w_0126_, w_0724_);
or (w_0777_, w_0741_, w_0549_);
or (w_0625_, w_0384_, w_0271_);
or (w_0676_, w_0093_, w_0582_);
not (w_0012_, w_0916_);
or (w_0065_, in15[4], w_0573_);
and (w_0539_, w_0447_, w_0419_);
or (w_0667_, w_0609_, w_0238_);
or (w_0843_, in12[5], w_0608_);
or (w_0837_, w_0839_, w_0326_);
and (w_0762_, in7[0], in8[0]);
not (w_0882_, w_0190_);
or (w_0460_, w_0467_, w_0883_);
or (w_0450_, w_0587_, w_0570_);
not (w_0572_, in11[3]);
and (w_0197_, w_0801_, w_0099_);
and (w_0438_, w_0126_, w_0724_);
and (w_0596_, w_0447_, w_0052_);
and (w_0405_, w_0904_, w_0072_);
or (w_0816_, w_0942_, w_0195_);
and (w_0616_, w_0206_, w_0026_);
or (w_0704_, w_0166_, w_0412_);
not (w_0440_, in12[3]);
and (w_0761_, w_0490_, w_0485_);
or (out12[0], w_0428_, w_0810_);
or (w_0305_, w_0015_, w_0284_);
and (w_0196_, in9[0], w_0123_);
or (w_0593_, w_0720_, w_0020_);
or (w_0944_, w_0349_, w_0824_);
or (w_0484_, w_0535_, w_0243_);
or (w_0296_, w_0509_, w_0307_);
and (w_0195_, w_0932_, w_0044_);
and (w_0629_, in13[1], in14[1]);
or (w_0442_, w_0074_, w_0768_);
and (w_0335_, w_0774_, w_0309_);
and (w_0509_, in15[3], w_0729_);
and (w_0823_, w_0169_, w_0372_);
not (w_0336_, w_0566_);
and (w_0371_, w_0525_, w_0670_);
and (w_0493_, w_0642_, w_0697_);
and (w_0885_, w_0852_, w_0843_);
and (w_0765_, w_0176_, w_0794_);
or (w_0604_, w_0884_, w_0792_);
and (w_0266_, w_0781_, w_0212_);
or (w_0419_, w_0567_, w_0047_);
and (w_0618_, w_0826_, w_0151_);
and (w_0430_, out4[0], w_0930_);
and (w_0734_, w_0051_, w_0367_);
not (w_0452_, in14[4]);
and (w_0949_, w_0893_, w_0898_);
and (w_0114_, w_0196_, w_0771_);
and (w_0186_, w_0239_, w_0530_);
and (w_0252_, in10[3], in11[3]);
and (w_0774_, w_0667_, w_0246_);
or (w_0767_, w_0837_, w_0004_);
not (w_0664_, w_0820_);
and (w_0889_, w_0504_, w_0784_);
or (w_0236_, w_0725_, w_0473_);
or (w_0844_, w_0000_, w_0744_);
and (w_0025_, w_0591_, w_0122_);
or (w_0627_, in9[2], w_0226_);
not (w_0225_, w_0201_);
and (w_0696_, w_0558_, w_0604_);
or (w_0630_, w_0869_, w_0227_);
not (w_0102_, w_0286_);
or (w_0640_, in3[2], w_0200_);
or (w_0673_, w_0011_, w_0106_);
or (w_0901_, w_0261_, w_0931_);
and (w_0459_, w_0444_, w_0730_);
or (w_0550_, w_0655_, w_0392_);
or (w_0660_, w_0869_, w_0538_);
and (w_0753_, w_0299_, w_0386_);
or (w_0112_, w_0412_, w_0085_);
and (w_0665_, w_0617_, w_0118_);
and (w_0522_, w_0415_, w_0071_);
and (w_0280_, w_0172_, w_0466_);
and (w_0850_, w_0813_, w_0783_);
and (w_0520_, w_0634_, w_0632_);
or (w_0510_, w_0224_, w_0515_);
not (w_0839_, in7[0]);
or (w_0289_, w_0770_, w_0139_);
or (w_0345_, w_0795_, w_0891_);
or (w_0904_, w_0357_, w_0914_);
not (w_0429_, w_0745_);
and (w_0738_, w_0088_, w_0393_);
or (w_0337_, w_0548_, w_0913_);
and (w_0538_, w_0716_, w_0554_);
and (w_0287_, w_0095_, w_0533_);
or (w_0921_, w_0400_, w_0125_);
and (w_0282_, w_0235_, w_0347_);
or (w_0678_, w_0059_, w_0800_);
or (w_0360_, w_0256_, w_0427_);
and (w_0498_, w_0306_, w_0510_);
and (w_0512_, w_0725_, w_0473_);
or (w_0019_, in12[3], w_0129_);
or (w_0570_, w_0196_, w_0228_);
or (w_0451_, in7[4], in8[4]);
and (w_0021_, w_0668_, w_0157_);
and (w_0022_, w_0248_, w_0694_);
not (w_0770_, in10[1]);
or (w_0913_, w_0430_, w_0511_);
or (w_0406_, w_0144_, w_0346_);
not (w_0836_, in7[1]);
or (w_0748_, w_0660_, w_0859_);
or (w_0383_, w_0305_, w_0132_);
or (w_0348_, w_0374_, w_0027_);
or (out12[2], w_0101_, w_0831_);
or (out13[0], w_0621_, w_0335_);
or (w_0216_, w_0908_, w_0665_);
not (w_0461_, w_0738_);
not (w_0387_, w_0939_);
not (w_0231_, w_0168_);
or (w_0127_, w_0791_, w_0303_);
and (w_0500_, w_0479_, w_0155_);
and (w_0927_, w_0135_, w_0623_);
not (w_0663_, w_0185_);
not (w_0699_, in3[1]);
and (w_0668_, w_0056_, w_0302_);
not (w_0087_, w_0749_);
or (w_0189_, w_0135_, w_0623_);
and (w_0215_, w_0109_, w_0445_);
and (w_0711_, w_0441_, w_0885_);
not (w_0242_, w_0305_);
not (w_0111_, w_0260_);
not (w_0390_, w_0119_);
or (w_0506_, in9[0], w_0123_);
not (w_0343_, w_0813_);
not (w_0792_, w_0527_);
and (w_0263_, w_0571_, w_0236_);
and (w_0899_, w_0051_, w_0474_);
and (w_0125_, w_0713_, w_0544_);
not (w_0852_, w_0535_);
or (w_0386_, w_0734_, w_0219_);
or (w_0652_, in7[0], in8[0]);
not (w_0851_, w_0499_);
or (w_0656_, w_0742_, w_0532_);
or (out8[0], w_0912_, w_0495_);
or (w_0353_, w_0077_, w_0508_);
or (w_0047_, w_0021_, w_0691_);
and (out11[2], w_0412_, w_0743_);
and (w_0448_, w_0689_, w_0638_);
not (w_0249_, w_0845_);
and (w_0691_, w_0234_, w_0469_);
or (w_0934_, w_0242_, w_0070_);
not (w_0329_, w_0455_);
or (w_0128_, w_0531_, w_0846_);
or (w_0780_, w_0261_, w_0409_);
not (w_0702_, in12[2]);
and (w_0175_, w_0797_, w_0487_);
and (w_0267_, w_0499_, w_0850_);
not (w_0074_, in15[6]);
or (w_0327_, in10[2], in11[2]);
and (w_0920_, in9[4], w_0943_);
and (w_0701_, w_0807_, w_0704_);
and (w_0511_, w_0551_, w_0045_);
or (w_0635_, w_0293_, w_0264_);
and (w_0626_, w_0593_, w_0752_);
or (w_0456_, w_0313_, w_0576_);
or (w_0281_, w_0774_, w_0309_);
and (w_0062_, in15[6], w_0266_);
or (w_0024_, in7[3], in8[3]);
and (w_0359_, w_0189_, w_0133_);
and (w_0395_, in10[1], in11[1]);
or (w_0801_, w_0198_, w_0208_);
and (w_0828_, w_0179_, w_0639_);
not (w_0004_, w_0643_);
not (w_0779_, w_0414_);
or (w_0818_, w_0183_, w_0494_);
or (w_0907_, w_0301_, w_0205_);
or (w_0815_, in13[0], in14[0]);
not (w_0726_, w_0188_);
and (w_0363_, w_0063_, w_0465_);
and (w_0183_, w_0893_, w_0866_);
not (w_0277_, w_0010_);
and (w_0575_, w_0153_, w_0454_);
and (w_0926_, w_0263_, w_0915_);
not (w_0113_, in14[1]);
or (w_0639_, w_0257_, w_0057_);
or (w_0122_, w_0270_, w_0498_);
and (w_0819_, in7[2], in8[2]);
or (w_0432_, w_0713_, w_0544_);
and (w_0445_, w_0801_, w_0076_);
or (w_0446_, w_0252_, w_0014_);
or (out3[1], w_0154_, w_0401_);
and (w_0130_, w_0807_, w_0595_);
not (w_0110_, w_0661_);
or (w_0870_, w_0463_, w_0856_);
and (w_0369_, w_0655_, w_0392_);
and (w_0607_, w_0328_, w_0832_);
or (w_0309_, w_0171_, w_0948_);
or (w_0536_, w_0306_, w_0510_);
not (w_0239_, w_0791_);
and (w_0079_, w_0407_, w_0677_);
not (w_0275_, in10[2]);
and (w_0653_, w_0616_, w_0073_);
and (w_0573_, w_0454_, w_0521_);
or (w_0425_, w_0916_, w_0114_);
and (w_0834_, w_0338_, w_0646_);
and (w_0166_, w_0551_, w_0683_);
or (w_0120_, w_0471_, w_0458_);
and (w_0162_, in15[5], w_0519_);
and (w_0613_, w_0571_, w_0797_);
and (w_0922_, w_0662_, w_0719_);
not (w_0407_, w_0059_);
and (w_0909_, w_0345_, w_0536_);
or (w_0308_, in13[5], in14[5]);
not (w_0918_, w_0934_);
and (w_0178_, w_0007_, w_0398_);
or (w_0617_, w_0941_, w_0542_);
or (w_0657_, w_0353_, w_0949_);
or (w_0712_, w_0802_, w_0277_);
or (w_0533_, w_0676_, w_0636_);
or (w_0291_, w_0426_, w_0193_);
or (w_0212_, w_0552_, w_0722_);
or (w_0477_, in4[1], in5[1]);
not (w_0674_, in5[2]);
or (w_0807_, w_0357_, w_0750_);
or (w_0404_, w_0875_, w_0351_);
or (w_0757_, w_0434_, w_0152_);
and (w_0716_, in4[0], in5[0]);
and (w_0144_, w_0216_, w_0006_);
or (w_0331_, w_0940_, w_0161_);
and (w_0006_, w_0793_, w_0829_);
or (w_0254_, w_0760_, w_0598_);
and (w_0086_, w_0300_, w_0686_);
and (w_0200_, w_0545_, w_0560_);
and (w_0067_, w_0820_, w_0303_);
and (w_0233_, out1[1], w_0028_);
or (w_0002_, in15[6], w_0266_);
and (w_0935_, w_0399_, w_0174_);
and (w_0027_, w_0345_, w_0379_);
or (w_0504_, w_0738_, w_0350_);
or (w_0039_, w_0400_, w_0505_);
or (w_0116_, in12[1], w_0010_);
and (w_0121_, w_0421_, w_0232_);
or (w_0623_, w_0688_, w_0923_);
not (w_0782_, w_0057_);
or (w_0878_, out1[1], w_0028_);
not (w_0295_, in15[4]);
or (w_0169_, w_0021_, w_0760_);
or (w_0155_, w_0276_, w_0756_);
not (w_0838_, in13[5]);
and (w_0464_, w_0787_, w_0529_);
and (w_0171_, w_0199_, w_0473_);
not (w_0013_, in11[4]);
and (w_0283_, w_0565_, w_0340_);
or (w_0560_, w_0635_, w_0079_);
and (w_0182_, w_0732_, w_0622_);
and (w_0097_, w_0574_, w_0001_);
not (w_0655_, in15[5]);
not (w_0811_, w_0648_);
and (w_0527_, w_0558_, w_0577_);
and (w_0190_, w_0620_, w_0425_);
or (w_0342_, w_0338_, w_0703_);
not (w_0937_, w_0840_);
or (w_0867_, w_0260_, w_0933_);
or (w_0525_, w_0897_, w_0375_);
and (w_0229_, w_0622_, w_0120_);
and (w_0115_, w_0772_, w_0815_);
and (w_0643_, w_0537_, w_0919_);
and (w_0368_, w_0726_, w_0009_);
and (w_0370_, w_0069_, w_0141_);
or (w_0561_, w_0039_, w_0922_);
and (w_0290_, w_0712_, w_0194_);
or (w_0421_, w_0772_, w_0365_);
or (out5[1], w_0754_, w_0083_);
and (w_0518_, w_0181_, w_0865_);
not (w_0515_, w_0379_);
and (w_0261_, w_0678_, w_0092_);
or (w_0788_, w_0803_, w_0382_);
or (w_0733_, w_0607_, w_0148_);
or (w_0133_, in15[2], w_0626_);
and (w_0000_, in15[0], w_0115_);
and (w_0156_, w_0261_, w_0931_);
not (w_0093_, in6[0]);
and (w_0766_, w_0419_, w_0054_);
not (w_0628_, w_0073_);
and (w_0492_, in12[1], w_0010_);
or (w_0785_, in3[0], w_0745_);
and (w_0585_, w_0557_, w_0041_);
or (w_0415_, w_0512_, w_0926_);
or (w_0165_, w_0166_, out1[1]);
and (w_0354_, w_0351_, w_0238_);
or (w_0812_, w_0616_, w_0234_);
not (w_0433_, w_0829_);
and (w_0848_, w_0100_, w_0896_);
not (w_0284_, w_0179_);
and (w_0203_, w_0107_, w_0405_);
or (w_0357_, out4[0], w_0333_);
or (w_0462_, in10[1], in11[1]);
and (w_0830_, w_0604_, w_0423_);
and (w_0742_, w_0289_, w_0938_);
not (w_0924_, in2[0]);
not (w_0056_, w_0711_);
or (w_0319_, w_0620_, w_0425_);
not (w_0507_, w_0041_);
or (w_0577_, in10[4], in11[4]);
and (w_0346_, w_0753_, w_0272_);
or (w_0080_, w_0088_, w_0393_);
or (w_0447_, w_0234_, w_0469_);
or (w_0092_, w_0741_, w_0438_);
or (w_0917_, w_0806_, w_0363_);
not (w_0063_, w_0819_);
or (w_0840_, in3[1], w_0464_);
and (w_0741_, in3[2], w_0200_);
or (w_0234_, w_0711_, w_0910_);
not (w_0070_, w_0132_);
not (w_0255_, w_0474_);
or (w_0141_, w_0043_, w_0259_);
or (w_0153_, w_0637_, w_0452_);
and (w_0247_, w_0552_, w_0722_);
and (w_0804_, w_0786_, w_0653_);
and (w_0351_, w_0780_, w_0334_);
or (w_0606_, w_0104_, w_0630_);
not (w_0005_, w_0391_);
and (w_0620_, w_0110_, w_0627_);
and (w_0720_, w_0574_, w_0421_);
or (w_0936_, w_0278_, w_0737_);
and (w_0916_, in9[1], w_0310_);
or (w_0862_, w_0177_, w_0899_);
or (w_0790_, w_0613_, w_0378_);
or (w_0473_, w_0516_, w_0553_);
not (w_0582_, w_0817_);
not (w_0434_, in4[1]);
and (w_0756_, w_0197_, w_0281_);
and (w_0517_, w_0036_, w_0576_);
or (w_0439_, w_0504_, w_0784_);
and (w_0729_, w_0536_, w_0348_);
and (w_0688_, w_0475_, w_0371_);
and (w_0090_, w_0229_, w_0366_);
not (w_0905_, w_0462_);
or (w_0095_, w_0269_, w_0779_);
and (w_0274_, in15[4], w_0573_);
or (w_0417_, w_0723_, w_0572_);
and (w_0103_, w_0295_, w_0798_);
not (w_0227_, w_0477_);
or (w_0362_, w_0929_, w_0134_);
or (w_0136_, in13[4], in14[4]);
and (w_0763_, w_0550_, w_0138_);
and (w_0603_, w_0575_, w_0871_);
or (w_0140_, w_0679_, w_0725_);
or (w_0915_, w_0381_, w_0814_);
or (w_0248_, w_0666_, w_0250_);
or (w_0752_, w_0475_, w_0371_);
or (w_0211_, w_0750_, w_0199_);
not (w_0841_, w_0701_);
and (w_0032_, w_0296_, w_0654_);
or (w_0638_, w_0575_, w_0871_);
or (w_0871_, w_0849_, w_0513_);
and (out11[1], w_0409_, w_0579_);
and (w_0942_, in15[1], w_0121_);
or (w_0041_, w_0813_, w_0783_);
and (w_0402_, w_0611_, w_0312_);
or (w_0046_, w_0685_, w_0736_);
or (out12[1], w_0067_, w_0180_);
or (w_0566_, w_0351_, w_0238_);
not (w_0778_, w_0754_);
and (w_0344_, w_0533_, w_0650_);
or (w_0551_, w_0342_, w_0754_);
or (w_0100_, w_0395_, w_0178_);
not (w_0089_, in12[4]);
or (w_0476_, w_0773_, w_0396_);
not (w_0037_, w_0783_);
or (w_0714_, w_0492_, w_0075_);
not (w_0903_, w_0147_);
or (w_0054_, w_0472_, w_0596_);
or (w_0602_, w_0936_, w_0182_);
and (w_0149_, w_0461_, w_0080_);
and (w_0377_, w_0662_, w_0586_);
and (w_0749_, w_0137_, out10[2]);
and (w_0401_, w_0347_, w_0684_);
and (w_0615_, w_0211_, w_0561_);
and (w_0449_, w_0201_, w_0853_);
or (w_0008_, in4[2], in5[2]);
or (w_0418_, w_0213_, w_0674_);
or (w_0044_, w_0035_, w_0081_);
or (w_0679_, w_0890_, w_0420_);
or (w_0670_, in13[2], in14[2]);
not (w_0322_, w_0015_);
not (w_0031_, in10[4]);
or (w_0559_, w_0137_, out10[2]);
or (w_0082_, w_0230_, w_0581_);
and (w_0771_, w_0012_, w_0017_);
and (w_0516_, w_0344_, w_0784_);
and (out7[1], w_0559_, w_0087_);
and (w_0469_, w_0682_, w_0119_);
or (w_0181_, w_0809_, w_0170_);
and (w_0592_, w_0870_, w_0667_);
or (w_0690_, w_0036_, w_0576_);
and (w_0600_, w_0418_, w_0360_);
and (w_0736_, w_0628_, w_0585_);
or (w_0241_, w_0705_, w_0924_);
and (w_0292_, w_0725_, w_0313_);
or (w_0523_, w_0942_, w_0739_);
and (w_0579_, w_0324_, w_0789_);
or (w_0060_, w_0548_, w_0766_);
or (w_0199_, w_0728_, w_0244_);
or (w_0358_, in10[5], in11[5]);
not (w_0933_, w_0669_);
or (w_0107_, w_0512_, w_0038_);
or (w_0396_, w_0188_, w_0633_);
or (w_0822_, w_0716_, w_0554_);
and (w_0416_, w_0613_, w_0378_);
and (w_0188_, in6[3], w_0709_);
not (w_0888_, w_0106_);
or (w_0893_, w_0591_, w_0122_);
and (w_0264_, w_0693_, w_0273_);
or (out2[1], w_0413_, w_0449_);
or (w_0257_, w_0819_, w_0648_);
and (w_0373_, in10[2], in11[2]);
and (w_0084_, in13[0], in14[0]);
or (w_0747_, w_0551_, w_0045_);
and (w_0154_, w_0050_, w_0042_);
and (w_0077_, in15[2], w_0626_);
or (w_0160_, w_0634_, w_0632_);
not (w_0549_, w_0640_);
and (w_0030_, w_0708_, w_0158_);
and (w_0073_, w_0499_, w_0265_);
and (w_0684_, w_0833_, w_0540_);
and (w_0278_, w_0279_, w_0601_);
or (w_0563_, in6[0], w_0817_);
or (w_0011_, w_0610_, w_0524_);
not (w_0723_, in10[3]);
or (w_0179_, w_0491_, w_0782_);
and (w_0276_, w_0879_, w_0867_);
not (w_0316_, w_0767_);
or (w_0503_, w_0355_, w_0820_);
and (w_0096_, w_0448_, w_0569_);
or (w_0033_, w_0699_, w_0502_);
and (out10[2], w_0561_, w_0432_);
or (w_0781_, w_0448_, w_0569_);
and (w_0361_, w_0360_, w_0748_);
and (w_0598_, w_0567_, w_0047_);
and (w_0259_, w_0679_, w_0583_);
and (w_0297_, w_0530_, w_0579_);
or (w_0177_, w_0492_, w_0834_);
and (w_0333_, w_0342_, w_0754_);
not (w_0703_, w_0697_);
or (w_0886_, w_0539_, w_0046_);
or (w_0845_, in6[1], w_0414_);
and (w_0148_, w_0731_, w_0769_);
or (w_0150_, w_0850_, w_0507_);
or (w_0001_, in13[1], in14[1]);
and (w_0118_, w_0299_, w_0019_);
and (w_0810_, w_0300_, w_0791_);
not (w_0750_, w_0412_);
and (w_0479_, w_0907_, w_0641_);
and (w_0007_, in10[0], in11[0]);
and (w_0881_, w_0794_, w_0788_);
not (w_0066_, w_0889_);
not (w_0833_, w_0114_);
not (w_0139_, in11[1]);
and (w_0746_, w_0676_, w_0636_);
and (w_0868_, w_0854_, w_0184_);
and (out9[1], w_0595_, w_0167_);
and (w_0035_, w_0084_, w_0097_);
or (w_0324_, w_0229_, w_0914_);
and (w_0634_, in3[0], w_0745_);
or (w_0051_, w_0702_, w_0005_);
not (w_0049_, w_0950_);
or (w_0017_, in9[1], w_0310_);
or (w_0708_, w_0645_, w_0777_);
or (w_0191_, w_0658_, w_0267_);
or (w_0544_, w_0349_, w_0325_);
or (w_0541_, w_0892_, w_0707_);
or (w_0020_, w_0675_, w_0078_);
or (w_0644_, w_0300_, w_0686_);
and (w_0524_, w_0446_, w_0527_);
and (w_0727_, w_0514_, w_0715_);
not (out4[0], w_0551_);
or (w_0485_, w_0332_, w_0763_);
and (w_0534_, w_0011_, w_0106_);
and (w_0576_, w_0695_, w_0160_);
and (w_0610_, in10[4], in11[4]);
not (w_0642_, w_0338_);
and (w_0508_, w_0523_, w_0359_);
and (w_0393_, w_0501_, w_0315_);
and (w_0293_, in1[1], in2[1]);
or (w_0557_, w_0343_, w_0037_);
or (out7[0], w_0173_, w_0117_);
and (w_0820_, w_0386_, w_0424_);
or (w_0185_, w_0535_, w_0711_);
and (w_0338_, in12[0], w_0590_);
and (w_0164_, w_0808_, w_0656_);
or (w_0945_, w_0415_, w_0071_);
and (w_0409_, w_0872_, w_0131_);
not (w_0221_, w_0368_);
or (w_0650_, w_0826_, w_0151_);
not (w_0721_, w_0686_);
and (w_0260_, w_0254_, w_0083_);
not (w_0427_, w_0859_);
or (w_0797_, w_0107_, w_0405_);
and (w_0306_, w_0525_, w_0593_);
or (w_0875_, w_0000_, w_0210_);
and (w_0101_, w_0279_, w_0355_);
and (w_0880_, w_0140_, w_0337_);
and (w_0068_, w_0237_, w_0016_);
and (w_0288_, w_0599_, w_0443_);
or (w_0094_, w_0209_, out1[0]);
and (w_0939_, in10[5], in11[5]);
and (w_0666_, w_0881_, w_0614_);
or (w_0474_, in12[2], w_0391_);
or (w_0376_, w_0426_, w_0145_);
or (w_0681_, w_0293_, w_0245_);
and (w_0724_, w_0411_, w_0640_);
or (w_0206_, w_0410_, w_0918_);
and (w_0391_, w_0656_, w_0671_);
or (w_0772_, w_0064_, w_0855_);
or (w_0340_, w_0162_, w_0369_);
and (w_0317_, w_0686_, w_0684_);
and (w_0381_, w_0166_, w_0706_);
not (w_0897_, in13[2]);
and (w_0632_, w_0033_, w_0840_);
and (w_0214_, w_0547_, w_0514_);
or (w_0706_, w_0233_, w_0517_);
and (w_0614_, w_0894_, w_0481_);
or (w_0584_, w_0600_, w_0877_);
or (w_0380_, in1[0], in2[0]);
not (w_0710_, in3[0]);
or (w_0299_, w_0440_, w_0740_);
and (w_0861_, w_0672_, w_0886_);
not (w_0078_, w_0670_);
or (w_0543_, w_0718_, w_0935_);
and (out11[0], w_0207_, w_0148_);
or (w_0172_, w_0162_, w_0285_);
and (w_0244_, w_0936_, w_0182_);
and (w_0739_, w_0000_, w_0744_);
and (w_0759_, out1[0], w_0928_);
and (w_0817_, w_0104_, w_0061_);
and (w_0658_, w_0851_, w_0557_);
and (w_0864_, in4[3], in5[3]);
or (w_0803_, w_0685_, w_0823_);
and (w_0486_, w_0456_, w_0946_);
and (w_0059_, in1[2], in2[2]);
or (w_0009_, in6[3], w_0709_);
or (w_0697_, in12[0], w_0590_);
or (w_0732_, w_0649_, w_0664_);
or (w_0798_, w_0068_, w_0578_);
not (w_0326_, in8[0]);
and (w_0645_, w_0033_, w_0695_);
or (w_0612_, w_0164_, w_0142_);
or (w_0157_, w_0280_, w_0390_);
not (w_0481_, w_0238_);
and (w_0180_, w_0664_, w_0530_);
and (w_0413_, w_0225_, w_0352_);
or (out5[0], w_0426_, w_0473_);
not (w_0633_, w_0872_);
and (w_0161_, w_0649_, w_0664_);
not (w_0855_, in14[0]);
and (w_0205_, w_0556_, w_0566_);
and (w_0578_, w_0909_, w_0082_);
or (w_0531_, w_0373_, w_0848_);
and (w_0554_, w_0757_, w_0477_);
or (w_0692_, w_0881_, w_0614_);
not (w_0857_, w_0019_);
or (w_0018_, w_0679_, w_0254_);
or (w_0641_, w_0248_, w_0694_);
or (w_0489_, w_0230_, w_0068_);
and (w_0014_, w_0531_, w_0846_);
and (w_0091_, w_0198_, w_0208_);
and (w_0713_, w_0211_, w_0112_);
and (w_0026_, w_0394_, w_0253_);
not (w_0799_, in13[1]);
or (w_0683_, w_0493_, w_0778_);
and (w_0431_, w_0651_, w_0298_);
or (w_0858_, in15[1], w_0121_);
and (w_0754_, w_0597_, w_0844_);
or (w_0698_, w_0661_, w_0190_);
and (w_0436_, w_0415_, w_0947_);
or (w_0872_, w_0217_, w_0221_);
or (w_0029_, w_0395_, w_0905_);
not (w_0556_, w_0354_);
and (w_0055_, w_0913_, w_0344_);
and (w_0279_, w_0589_, w_0262_);
and (w_0914_, w_0690_, w_0878_);
or (w_0789_, w_0181_, w_0706_);
or (w_0808_, w_0275_, w_0388_);
or (w_0842_, w_0932_, w_0044_);
and (w_0350_, w_0287_, w_0625_);
or (w_0076_, w_0925_, w_0621_);
or (w_0829_, in12[4], w_0830_);
or (w_0379_, in13[3], in14[3]);
or (w_0163_, w_0364_, w_0937_);
or (w_0540_, w_0196_, w_0771_);
or (out10[1], w_0156_, w_0108_);
or (out14[1], w_0804_, w_0329_);
and (w_0865_, w_0066_, w_0439_);
or (w_0443_, w_0086_, w_0430_);
or (w_0147_, in13[6], in14[6]);
or (w_0050_, w_0522_, w_0416_);
or (w_0392_, w_0496_, w_0603_);
or (w_0928_, w_0926_, w_0203_);
not (w_0064_, in13[0]);
and (w_0384_, in6[2], w_0361_);
or (w_0735_, w_0613_, w_0680_);
not (w_0375_, in14[2]);
and (w_0910_, w_0847_, w_0484_);
and (w_0414_, w_0606_, w_0822_);
not (w_0108_, w_0901_);
or (w_0237_, w_0224_, w_0270_);
or (w_0494_, w_0274_, w_0103_);
or (w_0787_, w_0241_, w_0681_);
and (w_0722_, w_0102_, w_0147_);
not (w_0042_, w_0684_);
or (out6[0], w_0403_, w_0385_);
and (w_0859_, w_0418_, w_0008_);
and (w_0887_, w_0645_, w_0777_);
and (w_0594_, w_0130_, w_0460_);
and (w_0755_, w_0168_, w_0528_);
not (w_0142_, w_0846_);
not (w_0929_, in1[1]);
or (w_0619_, w_0696_, w_0888_);
or (w_0894_, w_0647_, w_0202_);
or (w_0589_, w_0753_, w_0272_);
and (w_0463_, w_0803_, w_0382_);
not (w_0659_, w_0000_);
or (w_0586_, w_0351_, w_0229_);
not (out1[1], w_0036_);
and (w_0480_, in6[1], w_0414_);
and (w_0760_, w_0472_, w_0596_);
and (w_0495_, w_0607_, w_0148_);
and (w_0923_, w_0720_, w_0020_);
or (w_0911_, w_0870_, w_0667_);
and (w_0611_, w_0842_, w_0597_);
and (w_0398_, w_0289_, w_0462_);
not (w_0341_, w_0785_);
or (w_0472_, w_0278_, w_0728_);
and (w_0693_, in1[0], in2[0]);
and (w_0226_, w_0811_, w_0917_);
and (w_0467_, w_0548_, w_0913_);
and (w_0796_, w_0478_, w_0223_);
and (w_0207_, w_0882_, w_0319_);
or (w_0453_, w_0296_, w_0654_);
and (w_0132_, w_0314_, w_0451_);
buf (out14[2], 1'h1);
endmodule
