module new_sub_module1(
    input wire [6:0] new_in1,
    input wire [6:0] new_in13,
    input wire [6:0] new_in15,
    input wire [6:0] new_in5,
    input wire [6:0] new_in7,
    input wire [6:0] new_in8,
    input wire [6:0] new_in9,
    input wire [7:0] new_in14,
    input wire [7:0] new_in16,
    input wire [7:0] new_in2,
    input wire [7:0] new_in21,
    input wire [7:0] new_in22,
    input wire [7:0] new_in24,
    input wire [7:0] new_in3,
    input wire [7:0] new_in4,
    input wire [8:0] new_in10,
    input wire [8:0] new_in11,
    input wire [8:0] new_in12,
    input wire [8:0] new_in17,
    input wire [8:0] new_in18,
    input wire [8:0] new_in19,
    input wire [8:0] new_in20,
    input wire [8:0] new_in23,
    input wire [8:0] new_in6,
    output wire [4:0] new_out15,
    output wire [4:0] new_out2,
    output wire [4:0] new_out3,
    output wire [4:0] new_out6,
    output wire [4:0] new_out7,
    output wire [5:0] new_out1,
    output wire [5:0] new_out10,
    output wire [5:0] new_out14,
    output wire [5:0] new_out16,
    output wire [5:0] new_out4,
    output wire [5:0] new_out9,
    output wire [6:0] new_out11,
    output wire [6:0] new_out12,
    output wire [6:0] new_out13,
    output wire [6:0] new_out17,
    output wire [6:0] new_out18,
    output wire [6:0] new_out5,
    output wire [6:0] new_out8
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
wire w_0945_;
wire w_0946_;
wire w_0947_;
wire w_0948_;
wire w_0949_;
wire w_0950_;
wire w_0951_;
wire w_0952_;
wire w_0953_;
wire w_0954_;
wire w_0955_;
wire w_0956_;
wire w_0957_;
wire w_0958_;
wire w_0959_;
wire w_0960_;
wire w_0961_;
wire w_0962_;
wire w_0963_;
wire w_0964_;
wire w_0965_;
wire w_0966_;
wire w_0967_;
wire w_0968_;
wire w_0969_;
wire w_0970_;
wire w_0971_;
wire w_0972_;
wire w_0973_;
wire w_0974_;
wire w_0975_;
wire w_0976_;
wire w_0977_;
wire w_0978_;
wire w_0979_;
wire w_0980_;
wire w_0981_;
wire w_0982_;
wire w_0983_;
wire w_0984_;
wire w_0985_;
wire w_0986_;
wire w_0987_;
wire w_0988_;
wire w_0989_;
wire w_0990_;
wire w_0991_;
wire w_0992_;
wire w_0993_;
wire w_0994_;
wire w_0995_;
wire w_0996_;
wire w_0997_;
wire w_0998_;
wire w_0999_;
wire w_1000_;
wire w_1001_;
wire w_1002_;
wire w_1003_;
wire w_1004_;
wire w_1005_;
wire w_1006_;
wire w_1007_;
wire w_1008_;
wire w_1009_;
wire w_1010_;
wire w_1011_;
wire w_1012_;
wire w_1013_;
wire w_1014_;
wire w_1015_;
wire w_1016_;
wire w_1017_;
wire w_1018_;
wire w_1019_;
wire w_1020_;
wire w_1021_;
wire w_1022_;
wire w_1023_;
wire w_1024_;
wire w_1025_;
wire w_1026_;
wire w_1027_;
wire w_1028_;
wire w_1029_;
wire w_1030_;
wire w_1031_;
wire w_1032_;
wire w_1033_;
wire w_1034_;
wire w_1035_;
wire w_1036_;
wire w_1037_;
wire w_1038_;
wire w_1039_;
wire w_1040_;
wire w_1041_;
wire w_1042_;
wire w_1043_;
wire w_1044_;
wire w_1045_;
wire w_1046_;
wire w_1047_;
wire w_1048_;
wire w_1049_;
wire w_1050_;
wire w_1051_;
wire w_1052_;
wire w_1053_;
wire w_1054_;
wire w_1055_;
wire w_1056_;
wire w_1057_;
wire w_1058_;
wire w_1059_;
wire w_1060_;
wire w_1061_;
wire w_1062_;
wire w_1063_;
wire w_1064_;
wire w_1065_;
wire w_1066_;
wire w_1067_;
wire w_1068_;
wire w_1069_;
wire w_1070_;
wire w_1071_;
wire w_1072_;
wire w_1073_;
wire w_1074_;
wire w_1075_;
wire w_1076_;
wire w_1077_;
wire w_1078_;
wire w_1079_;
wire w_1080_;
wire w_1081_;
wire w_1082_;
wire w_1083_;
wire w_1084_;
wire w_1085_;
wire w_1086_;
wire w_1087_;
wire w_1088_;
wire w_1089_;
wire w_1090_;
wire w_1091_;
wire w_1092_;
wire w_1093_;
wire w_1094_;
wire w_1095_;
wire w_1096_;
wire w_1097_;
wire w_1098_;
wire w_1099_;
wire w_1100_;
wire w_1101_;
wire w_1102_;
wire w_1103_;
wire w_1104_;
wire w_1105_;
wire w_1106_;
wire w_1107_;
wire w_1108_;
wire w_1109_;
wire w_1110_;
wire w_1111_;
wire w_1112_;
wire w_1113_;
wire w_1114_;
wire w_1115_;
wire w_1116_;
wire w_1117_;
wire w_1118_;
wire w_1119_;
wire w_1120_;
wire w_1121_;
wire w_1122_;
wire w_1123_;
wire w_1124_;
wire w_1125_;
wire w_1126_;
wire w_1127_;
wire w_1128_;
wire w_1129_;
wire w_1130_;
wire w_1131_;
wire w_1132_;
wire w_1133_;
wire w_1134_;
wire w_1135_;
wire w_1136_;
wire w_1137_;
wire w_1138_;
wire w_1139_;
wire w_1140_;
wire w_1141_;
wire w_1142_;
wire w_1143_;
wire w_1144_;
wire w_1145_;
wire w_1146_;
wire w_1147_;
wire w_1148_;
wire w_1149_;
wire w_1150_;
wire w_1151_;
wire w_1152_;
wire w_1153_;
wire w_1154_;
wire w_1155_;
wire w_1156_;
wire w_1157_;
wire w_1158_;
wire w_1159_;
wire w_1160_;
wire w_1161_;
wire w_1162_;
wire w_1163_;
wire w_1164_;
wire w_1165_;
wire w_1166_;
wire w_1167_;
wire w_1168_;
wire w_1169_;
wire w_1170_;
wire w_1171_;
wire w_1172_;
wire w_1173_;
wire w_1174_;
wire w_1175_;
wire w_1176_;
wire w_1177_;
wire w_1178_;
wire w_1179_;
wire w_1180_;
wire w_1181_;
wire w_1182_;
wire w_1183_;
wire w_1184_;
wire w_1185_;
wire w_1186_;
wire w_1187_;
wire w_1188_;
wire w_1189_;
wire w_1190_;
wire w_1191_;
wire w_1192_;
wire w_1193_;
wire w_1194_;
wire w_1195_;
wire w_1196_;
wire w_1197_;
wire w_1198_;
wire w_1199_;
wire w_1200_;
wire w_1201_;
wire w_1202_;
wire w_1203_;
wire w_1204_;
wire w_1205_;
wire w_1206_;
wire w_1207_;
wire w_1208_;
wire w_1209_;
wire w_1210_;
wire w_1211_;
wire w_1212_;
wire w_1213_;
wire w_1214_;
wire w_1215_;
wire w_1216_;
wire w_1217_;
wire w_1218_;
wire w_1219_;
wire w_1220_;
wire w_1221_;
wire w_1222_;
wire w_1223_;
wire w_1224_;
wire w_1225_;
wire w_1226_;
wire w_1227_;
wire w_1228_;
wire w_1229_;
wire w_1230_;
wire w_1231_;
wire w_1232_;
wire w_1233_;
wire w_1234_;
wire w_1235_;
wire w_1236_;
wire w_1237_;
wire w_1238_;
wire w_1239_;
wire w_1240_;
wire w_1241_;
wire w_1242_;
wire w_1243_;
wire w_1244_;
wire w_1245_;
wire w_1246_;
wire w_1247_;
wire w_1248_;
wire w_1249_;
wire w_1250_;
wire w_1251_;
wire w_1252_;
wire w_1253_;
wire w_1254_;
wire w_1255_;
wire w_1256_;
wire w_1257_;
wire w_1258_;
wire w_1259_;
wire w_1260_;
wire w_1261_;
wire w_1262_;
wire w_1263_;
wire w_1264_;
wire w_1265_;
wire w_1266_;
wire w_1267_;
wire w_1268_;
wire w_1269_;
wire w_1270_;
wire w_1271_;
wire w_1272_;
wire w_1273_;
wire w_1274_;
wire w_1275_;
wire w_1276_;
wire w_1277_;
wire w_1278_;
wire w_1279_;
wire w_1280_;
wire w_1281_;
wire w_1282_;
wire w_1283_;
wire w_1284_;
wire w_1285_;
wire w_1286_;
wire w_1287_;
wire w_1288_;
wire w_1289_;
wire w_1290_;
wire w_1291_;
wire w_1292_;
wire w_1293_;
wire w_1294_;
wire w_1295_;
wire w_1296_;
wire w_1297_;
wire w_1298_;
wire w_1299_;
wire w_1300_;
wire w_1301_;
wire w_1302_;
wire w_1303_;
wire w_1304_;
wire w_1305_;
wire w_1306_;
wire w_1307_;
wire w_1308_;
wire w_1309_;
wire w_1310_;
wire w_1311_;
wire w_1312_;
wire w_1313_;
wire w_1314_;
wire w_1315_;
wire w_1316_;
wire w_1317_;
wire w_1318_;
wire w_1319_;
wire w_1320_;
wire w_1321_;
wire w_1322_;
wire w_1323_;
wire w_1324_;
wire w_1325_;
wire w_1326_;
wire w_1327_;
wire w_1328_;
wire w_1329_;
wire w_1330_;
wire w_1331_;
wire w_1332_;
wire w_1333_;
wire w_1334_;
wire w_1335_;
wire w_1336_;
wire w_1337_;
wire w_1338_;
wire w_1339_;
wire w_1340_;
wire w_1341_;
wire w_1342_;
wire w_1343_;
wire w_1344_;
wire w_1345_;
wire w_1346_;
wire w_1347_;
wire w_1348_;
wire w_1349_;
wire w_1350_;
wire w_1351_;
wire w_1352_;
wire w_1353_;
wire w_1354_;
wire w_1355_;
wire w_1356_;
wire w_1357_;
wire w_1358_;
wire w_1359_;
wire w_1360_;
wire w_1361_;
wire w_1362_;
wire w_1363_;
wire w_1364_;
wire w_1365_;
wire w_1366_;
wire w_1367_;
wire w_1368_;
wire w_1369_;
wire w_1370_;
wire w_1371_;
wire w_1372_;
wire w_1373_;
wire w_1374_;
wire w_1375_;
wire w_1376_;
wire w_1377_;
wire w_1378_;
wire w_1379_;
wire w_1380_;
wire w_1381_;
wire w_1382_;
wire w_1383_;
wire w_1384_;
wire w_1385_;
wire w_1386_;
wire w_1387_;
wire w_1388_;
wire w_1389_;
wire w_1390_;
wire w_1391_;
wire w_1392_;
wire w_1393_;
wire w_1394_;
wire w_1395_;
wire w_1396_;
wire w_1397_;
wire w_1398_;
wire w_1399_;
wire w_1400_;
wire w_1401_;
wire w_1402_;
wire w_1403_;
wire w_1404_;
wire w_1405_;
wire w_1406_;
wire w_1407_;
wire w_1408_;
wire w_1409_;
wire w_1410_;
wire w_1411_;
wire w_1412_;
wire w_1413_;
wire w_1414_;
wire w_1415_;
wire w_1416_;
wire w_1417_;
wire w_1418_;
wire w_1419_;
wire w_1420_;
wire w_1421_;
wire w_1422_;
wire w_1423_;
wire w_1424_;
wire w_1425_;
wire w_1426_;
wire w_1427_;
wire w_1428_;
wire w_1429_;
wire w_1430_;
wire w_1431_;
wire w_1432_;
wire w_1433_;
wire w_1434_;
wire w_1435_;
wire w_1436_;
wire w_1437_;
wire w_1438_;
wire w_1439_;
wire w_1440_;
wire w_1441_;
wire w_1442_;
wire w_1443_;
wire w_1444_;
wire w_1445_;
wire w_1446_;
wire w_1447_;
wire w_1448_;
wire w_1449_;
wire w_1450_;
wire w_1451_;
wire w_1452_;
wire w_1453_;
wire w_1454_;
wire w_1455_;
wire w_1456_;
wire w_1457_;
wire w_1458_;
wire w_1459_;
wire w_1460_;
wire w_1461_;
wire w_1462_;
wire w_1463_;
wire w_1464_;
wire w_1465_;
wire w_1466_;
wire w_1467_;
wire w_1468_;
wire w_1469_;
wire w_1470_;
wire w_1471_;
wire w_1472_;
wire w_1473_;
wire w_1474_;
wire w_1475_;
wire w_1476_;
wire w_1477_;
wire w_1478_;
wire w_1479_;
wire w_1480_;
wire w_1481_;
wire w_1482_;
wire w_1483_;
wire w_1484_;
wire w_1485_;
wire w_1486_;
wire w_1487_;
wire w_1488_;
wire w_1489_;
wire w_1490_;
wire w_1491_;
wire w_1492_;
wire w_1493_;
wire w_1494_;
wire w_1495_;
wire w_1496_;
wire w_1497_;
wire w_1498_;
wire w_1499_;
wire w_1500_;
wire w_1501_;
wire w_1502_;
wire w_1503_;
wire w_1504_;
wire w_1505_;
wire w_1506_;
wire w_1507_;
wire w_1508_;
wire w_1509_;
wire w_1510_;
wire w_1511_;
wire w_1512_;
wire w_1513_;
wire w_1514_;
wire w_1515_;
wire w_1516_;
wire w_1517_;
wire w_1518_;
wire w_1519_;
wire w_1520_;
wire w_1521_;
wire w_1522_;
wire w_1523_;
wire w_1524_;
wire w_1525_;
wire w_1526_;
wire w_1527_;
wire w_1528_;
wire w_1529_;
wire w_1530_;
wire w_1531_;
wire w_1532_;
wire w_1533_;
wire w_1534_;
wire w_1535_;
wire w_1536_;
wire w_1537_;
wire w_1538_;
wire w_1539_;
wire w_1540_;
wire w_1541_;
wire w_1542_;
wire w_1543_;
wire w_1544_;
wire w_1545_;
wire w_1546_;
wire w_1547_;
wire w_1548_;
wire w_1549_;
wire w_1550_;
wire w_1551_;
wire w_1552_;
wire w_1553_;
wire w_1554_;
wire w_1555_;
wire w_1556_;
wire w_1557_;
wire w_1558_;
wire w_1559_;
wire w_1560_;
wire w_1561_;
wire w_1562_;
wire w_1563_;
wire w_1564_;
wire w_1565_;
wire w_1566_;
wire w_1567_;
wire w_1568_;
wire w_1569_;
wire w_1570_;
wire w_1571_;
wire w_1572_;
wire w_1573_;
wire w_1574_;
wire w_1575_;
wire w_1576_;
wire w_1577_;
wire w_1578_;
wire w_1579_;
wire w_1580_;
wire w_1581_;
wire w_1582_;
wire w_1583_;
wire w_1584_;
wire w_1585_;
wire w_1586_;
wire w_1587_;
wire w_1588_;
wire w_1589_;
wire w_1590_;
wire w_1591_;
wire w_1592_;
wire w_1593_;
wire w_1594_;
wire w_1595_;
wire w_1596_;
wire w_1597_;
wire w_1598_;
wire w_1599_;
wire w_1600_;
wire w_1601_;
wire w_1602_;
wire w_1603_;
wire w_1604_;
wire w_1605_;
wire w_1606_;
wire w_1607_;
wire w_1608_;
wire w_1609_;
wire w_1610_;
wire w_1611_;
wire w_1612_;
wire w_1613_;
wire w_1614_;
wire w_1615_;
wire w_1616_;
wire w_1617_;
wire w_1618_;
wire w_1619_;
wire w_1620_;
wire w_1621_;
wire w_1622_;
wire w_1623_;
wire w_1624_;
wire w_1625_;
wire w_1626_;
wire w_1627_;
wire w_1628_;
wire w_1629_;
wire w_1630_;
wire w_1631_;
wire w_1632_;
wire w_1633_;
wire w_1634_;
wire w_1635_;
wire w_1636_;
wire w_1637_;
wire w_1638_;
wire w_1639_;
wire w_1640_;
wire w_1641_;
wire w_1642_;
wire w_1643_;
wire w_1644_;
wire w_1645_;
wire w_1646_;
wire w_1647_;
wire w_1648_;
wire w_1649_;
wire w_1650_;
wire w_1651_;
wire w_1652_;
wire w_1653_;
wire w_1654_;
wire w_1655_;
wire w_1656_;
wire w_1657_;
wire w_1658_;
wire w_1659_;
wire w_1660_;
wire w_1661_;
wire w_1662_;
wire w_1663_;
wire w_1664_;
wire w_1665_;
wire w_1666_;
wire w_1667_;
wire w_1668_;
wire w_1669_;
wire w_1670_;
wire w_1671_;
wire w_1672_;
wire w_1673_;
wire w_1674_;
wire w_1675_;
wire w_1676_;
wire w_1677_;
wire w_1678_;
wire w_1679_;
wire w_1680_;
wire w_1681_;
wire w_1682_;
wire w_1683_;
wire w_1684_;
wire w_1685_;
wire w_1686_;
wire w_1687_;
wire w_1688_;
wire w_1689_;
wire w_1690_;
wire w_1691_;
wire w_1692_;
wire w_1693_;
wire w_1694_;
wire w_1695_;
wire w_1696_;
wire w_1697_;
wire w_1698_;
wire w_1699_;
wire w_1700_;
wire w_1701_;
wire w_1702_;
wire w_1703_;
wire w_1704_;
wire w_1705_;
wire w_1706_;
wire w_1707_;
wire w_1708_;
wire w_1709_;
wire w_1710_;
wire w_1711_;
wire w_1712_;
wire w_1713_;
wire w_1714_;
wire w_1715_;
wire w_1716_;
wire w_1717_;
wire w_1718_;
wire w_1719_;
wire w_1720_;
wire w_1721_;
wire w_1722_;
wire w_1723_;
wire w_1724_;
wire w_1725_;
wire w_1726_;
wire w_1727_;
wire w_1728_;
wire w_1729_;
wire w_1730_;
wire w_1731_;
wire w_1732_;
wire w_1733_;
wire w_1734_;
wire w_1735_;
wire w_1736_;
wire w_1737_;
wire w_1738_;
wire w_1739_;
wire w_1740_;
wire w_1741_;
wire w_1742_;
wire w_1743_;
wire w_1744_;
wire w_1745_;
wire w_1746_;
wire w_1747_;
wire w_1748_;
wire w_1749_;
wire w_1750_;
wire w_1751_;
wire w_1752_;
wire w_1753_;
wire w_1754_;
wire w_1755_;
wire w_1756_;
wire w_1757_;
wire w_1758_;
wire w_1759_;
wire w_1760_;
wire w_1761_;
wire w_1762_;
wire w_1763_;
wire w_1764_;
wire w_1765_;
wire w_1766_;
wire w_1767_;
wire w_1768_;
wire w_1769_;
wire w_1770_;
wire w_1771_;
wire w_1772_;
wire w_1773_;
wire w_1774_;
wire w_1775_;
wire w_1776_;
wire w_1777_;
wire w_1778_;
wire w_1779_;
wire w_1780_;
wire w_1781_;
wire w_1782_;
wire w_1783_;
wire w_1784_;
wire w_1785_;
wire w_1786_;
wire w_1787_;
wire w_1788_;
wire w_1789_;
wire w_1790_;
wire w_1791_;
wire w_1792_;
wire w_1793_;
wire w_1794_;
wire w_1795_;
wire w_1796_;
wire w_1797_;
wire w_1798_;
wire w_1799_;
wire w_1800_;
wire w_1801_;
wire w_1802_;
wire w_1803_;
wire w_1804_;
wire w_1805_;
wire w_1806_;
wire w_1807_;
wire w_1808_;
wire w_1809_;
wire w_1810_;
wire w_1811_;
wire w_1812_;
wire w_1813_;
wire w_1814_;
wire w_1815_;
wire w_1816_;
wire w_1817_;
wire w_1818_;
wire w_1819_;
wire w_1820_;
wire w_1821_;
wire w_1822_;
wire w_1823_;
wire w_1824_;
wire w_1825_;
wire w_1826_;
wire w_1827_;
wire w_1828_;
wire w_1829_;
wire w_1830_;
wire w_1831_;
wire w_1832_;
wire w_1833_;
wire w_1834_;
wire w_1835_;
wire w_1836_;
wire w_1837_;
wire w_1838_;
wire w_1839_;
wire w_1840_;
wire w_1841_;
wire w_1842_;
wire w_1843_;
wire w_1844_;
wire w_1845_;
wire w_1846_;
wire w_1847_;
wire w_1848_;
wire w_1849_;
wire w_1850_;
wire w_1851_;
wire w_1852_;
wire w_1853_;
wire w_1854_;
wire w_1855_;
wire w_1856_;
wire w_1857_;
wire w_1858_;
wire w_1859_;
wire w_1860_;
wire w_1861_;
wire w_1862_;
wire w_1863_;
wire w_1864_;
wire w_1865_;
wire w_1866_;
wire w_1867_;
wire w_1868_;
wire w_1869_;
wire w_1870_;
wire w_1871_;
wire w_1872_;
wire w_1873_;
wire w_1874_;
wire w_1875_;
wire w_1876_;
wire w_1877_;
wire w_1878_;
wire w_1879_;
wire w_1880_;
wire w_1881_;
wire w_1882_;
wire w_1883_;
wire w_1884_;
wire w_1885_;
wire w_1886_;
wire w_1887_;
wire w_1888_;
wire w_1889_;
wire w_1890_;
wire w_1891_;
wire w_1892_;
wire w_1893_;
wire w_1894_;
wire w_1895_;
wire w_1896_;
wire w_1897_;
wire w_1898_;
wire w_1899_;
wire w_1900_;
wire w_1901_;
wire w_1902_;
wire w_1903_;
wire w_1904_;
wire w_1905_;
wire w_1906_;
wire w_1907_;
wire w_1908_;
wire w_1909_;
wire w_1910_;
wire w_1911_;
wire w_1912_;
wire w_1913_;
wire w_1914_;
wire w_1915_;
wire w_1916_;
wire w_1917_;
wire w_1918_;
wire w_1919_;
wire w_1920_;
wire w_1921_;
wire w_1922_;
wire w_1923_;
wire w_1924_;
wire w_1925_;
wire w_1926_;
wire w_1927_;
wire w_1928_;
wire w_1929_;
wire w_1930_;
wire w_1931_;
wire w_1932_;
wire w_1933_;
wire w_1934_;
wire w_1935_;
wire w_1936_;
wire w_1937_;
wire w_1938_;
wire w_1939_;
wire w_1940_;
wire w_1941_;
wire w_1942_;
wire w_1943_;
wire w_1944_;
wire w_1945_;
wire w_1946_;
wire w_1947_;
wire w_1948_;
wire w_1949_;
wire w_1950_;
wire w_1951_;
wire w_1952_;
wire w_1953_;
wire w_1954_;
wire w_1955_;
wire w_1956_;
wire w_1957_;
wire w_1958_;
wire w_1959_;
wire w_1960_;
wire w_1961_;
wire w_1962_;
wire w_1963_;
wire w_1964_;
wire w_1965_;
wire w_1966_;
wire w_1967_;
wire w_1968_;
wire w_1969_;
wire w_1970_;
wire w_1971_;
wire w_1972_;
wire w_1973_;
wire w_1974_;
wire w_1975_;
wire w_1976_;
wire w_1977_;
wire w_1978_;
wire w_1979_;
wire w_1980_;
wire w_1981_;
wire w_1982_;
wire w_1983_;
wire w_1984_;
wire w_1985_;
wire w_1986_;
wire w_1987_;
wire w_1988_;
wire w_1989_;
wire w_1990_;
wire w_1991_;
wire w_1992_;
wire w_1993_;
wire w_1994_;
wire w_1995_;
wire w_1996_;
wire w_1997_;
wire w_1998_;
wire w_1999_;
wire w_2000_;
wire w_2001_;
wire w_2002_;
wire w_2003_;
wire w_2004_;
wire w_2005_;
wire w_2006_;
wire w_2007_;
wire w_2008_;
wire w_2009_;
wire w_2010_;
wire w_2011_;
wire w_2012_;
wire w_2013_;
wire w_2014_;
wire w_2015_;
wire w_2016_;
wire w_2017_;
wire w_2018_;
wire w_2019_;
wire w_2020_;
wire w_2021_;
wire w_2022_;
wire w_2023_;
wire w_2024_;
wire w_2025_;
wire w_2026_;
wire w_2027_;
wire w_2028_;
wire w_2029_;
wire w_2030_;
wire w_2031_;
wire w_2032_;
wire w_2033_;
wire w_2034_;
wire w_2035_;
wire w_2036_;
wire w_2037_;
wire w_2038_;
wire w_2039_;
wire w_2040_;
wire w_2041_;
wire w_2042_;
wire w_2043_;
wire w_2044_;
wire w_2045_;
wire w_2046_;
wire w_2047_;
wire w_2048_;
wire w_2049_;
wire w_2050_;
wire w_2051_;
wire w_2052_;
wire w_2053_;
wire w_2054_;
wire w_2055_;
wire w_2056_;
wire w_2057_;
wire w_2058_;
wire w_2059_;
wire w_2060_;
wire w_2061_;
wire w_2062_;
wire w_2063_;
wire w_2064_;
wire w_2065_;
wire w_2066_;
wire w_2067_;
wire w_2068_;
wire w_2069_;
wire w_2070_;
wire w_2071_;
wire w_2072_;
wire w_2073_;
wire w_2074_;
wire w_2075_;
wire w_2076_;
wire w_2077_;
wire w_2078_;
wire w_2079_;
wire w_2080_;
wire w_2081_;
wire w_2082_;
wire w_2083_;
wire w_2084_;
wire w_2085_;
wire w_2086_;
wire w_2087_;
wire w_2088_;
wire w_2089_;
wire w_2090_;
wire w_2091_;
wire w_2092_;
wire w_2093_;
wire w_2094_;
wire w_2095_;
wire w_2096_;
wire w_2097_;
wire w_2098_;
wire w_2099_;
wire w_2100_;
wire w_2101_;
wire w_2102_;
wire w_2103_;
wire w_2104_;
wire w_2105_;
wire w_2106_;
wire w_2107_;
wire w_2108_;
wire w_2109_;
wire w_2110_;
wire w_2111_;
wire w_2112_;
wire w_2113_;
wire w_2114_;
wire w_2115_;
wire w_2116_;
wire w_2117_;
wire w_2118_;
wire w_2119_;
wire w_2120_;
wire w_2121_;
wire w_2122_;
wire w_2123_;
wire w_2124_;
wire w_2125_;
wire w_2126_;
wire w_2127_;
wire w_2128_;
wire w_2129_;
wire w_2130_;
wire w_2131_;
wire w_2132_;
wire w_2133_;
wire w_2134_;
wire w_2135_;
wire w_2136_;
wire w_2137_;
wire w_2138_;
wire w_2139_;
wire w_2140_;
wire w_2141_;
wire w_2142_;
wire w_2143_;
wire w_2144_;
wire w_2145_;
wire w_2146_;
wire w_2147_;
wire w_2148_;
wire w_2149_;
wire w_2150_;
wire w_2151_;
wire w_2152_;
wire w_2153_;
wire w_2154_;
wire w_2155_;
wire w_2156_;
wire w_2157_;
wire w_2158_;
wire w_2159_;
wire w_2160_;
wire w_2161_;
wire w_2162_;
wire w_2163_;
wire w_2164_;
wire w_2165_;
wire w_2166_;
wire w_2167_;
wire w_2168_;
wire w_2169_;
wire w_2170_;
wire w_2171_;
wire w_2172_;
wire w_2173_;
wire w_2174_;
wire w_2175_;
wire w_2176_;
wire w_2177_;
wire w_2178_;
wire w_2179_;
wire w_2180_;
wire w_2181_;
wire w_2182_;
wire w_2183_;
wire w_2184_;
wire w_2185_;
wire w_2186_;
wire w_2187_;
wire w_2188_;
wire w_2189_;
wire w_2190_;
wire w_2191_;
wire w_2192_;
wire w_2193_;
wire w_2194_;
wire w_2195_;
wire w_2196_;
wire w_2197_;
wire w_2198_;
wire w_2199_;
wire w_2200_;
wire w_2201_;
wire w_2202_;
wire w_2203_;
wire w_2204_;
wire w_2205_;
wire w_2206_;
wire w_2207_;
wire w_2208_;
wire w_2209_;
wire w_2210_;
wire w_2211_;
wire w_2212_;
wire w_2213_;
wire w_2214_;
wire w_2215_;
wire w_2216_;
wire w_2217_;
wire w_2218_;
wire w_2219_;
wire w_2220_;
wire w_2221_;
wire w_2222_;
wire w_2223_;
wire w_2224_;
wire w_2225_;
wire w_2226_;
wire w_2227_;
wire w_2228_;
wire w_2229_;
wire w_2230_;
wire w_2231_;
wire w_2232_;
wire w_2233_;
wire w_2234_;
wire w_2235_;
wire w_2236_;
wire w_2237_;
wire w_2238_;
wire w_2239_;
wire w_2240_;
wire w_2241_;
wire w_2242_;
wire w_2243_;
wire w_2244_;
wire w_2245_;
wire w_2246_;
wire w_2247_;
wire w_2248_;
wire w_2249_;
wire w_2250_;
wire w_2251_;
wire w_2252_;
wire w_2253_;
wire w_2254_;
wire w_2255_;
wire w_2256_;
wire w_2257_;
wire w_2258_;
wire w_2259_;
wire w_2260_;
wire w_2261_;
wire w_2262_;
wire w_2263_;
wire w_2264_;
wire w_2265_;
wire w_2266_;
wire w_2267_;
wire w_2268_;
wire w_2269_;
wire w_2270_;
wire w_2271_;
wire w_2272_;
wire w_2273_;
wire w_2274_;
wire w_2275_;
wire w_2276_;
wire w_2277_;
wire w_2278_;
wire w_2279_;
wire w_2280_;
wire w_2281_;
wire w_2282_;
wire w_2283_;
wire w_2284_;
wire w_2285_;
wire w_2286_;
wire w_2287_;
wire w_2288_;
wire w_2289_;
wire w_2290_;
wire w_2291_;
wire w_2292_;
wire w_2293_;
wire w_2294_;
wire w_2295_;
wire w_2296_;
wire w_2297_;
wire w_2298_;
wire w_2299_;
wire w_2300_;
wire w_2301_;
wire w_2302_;
wire w_2303_;
wire w_2304_;
wire w_2305_;
wire w_2306_;
wire w_2307_;
wire w_2308_;
wire w_2309_;
wire w_2310_;
wire w_2311_;
wire w_2312_;
wire w_2313_;
wire w_2314_;
wire w_2315_;
wire w_2316_;
wire w_2317_;
wire w_2318_;
wire w_2319_;
wire w_2320_;
wire w_2321_;
wire w_2322_;
wire w_2323_;
wire w_2324_;
or (w_1195_, new_in22[0], new_in16[0]);
nand (w_1179_, new_in16[7], w_0705_);
xor (w_0444_, new_in11[2], w_0785_);
nand (w_0518_, w_0808_, w_0551_);
not (w_0321_, w_1368_);
and (w_0122_, w_0003_, w_0859_);
nand (w_0131_, new_in23[4], new_in6[4]);
and (w_0319_, w_0531_, w_0082_);
xor (w_1557_, w_1846_, w_1010_);
nand (w_0177_, w_1905_, w_0288_);
nand (w_1246_, w_0825_, w_1498_);
nand (w_1322_, new_in10[8], w_0434_);
or (w_1294_, w_0789_, w_1913_);
nand (w_0336_, w_1528_, w_1948_);
and (w_0503_, new_in5[6], w_1200_);
nand (w_0273_, w_0997_, w_1197_);
nand (w_1450_, w_1784_, w_0786_);
and (new_out8[3], w_1976_, w_1096_);
nand (w_0068_, w_1234_, w_0252_);
nand (w_1953_, new_in16[7], w_0860_);
nand (w_0089_, w_1499_, w_0684_);
xor (w_1616_, new_in19[2], new_in6[1]);
and (w_1632_, w_1234_, w_0662_);
or (w_1664_, new_in21[0], w_1960_);
nand (new_out13[2], w_1501_, w_1341_);
and (w_1771_, new_in16[7], w_2250_);
nand (w_0402_, new_in22[5], new_in9[2]);
and (w_2313_, w_1203_, w_1094_);
and (w_0338_, w_2124_, w_0155_);
and (w_1905_, new_in10[8], w_1231_);
nand (w_1502_, w_0680_, w_1559_);
and (new_out2[3], w_0624_, w_1610_);
and (w_1680_, w_0132_, w_0704_);
xor (w_2063_, new_in23[3], new_in12[3]);
nand (w_0255_, w_0558_, w_1393_);
nand (w_0378_, w_0890_, w_0236_);
xor (w_1560_, w_1995_, w_1987_);
xor (w_0605_, w_1211_, w_0040_);
and (w_0759_, w_0338_, w_0480_);
and (w_1062_, new_in5[6], w_1382_);
nor (new_out5[3], w_1603_, w_1651_);
or (w_0890_, w_0263_, w_1522_);
nand (w_1665_, w_0602_, w_0538_);
nand (w_1336_, new_in13[4], new_in1[4]);
and (w_0384_, w_2121_, w_0751_);
or (w_0886_, w_2114_, w_2126_);
xor (w_0970_, w_1441_, w_0546_);
and (w_1024_, w_2093_, w_0234_);
nand (w_0813_, w_1231_, w_0617_);
and (w_0806_, new_in5[3], w_1695_);
nand (w_0433_, w_0738_, w_1697_);
and (w_0330_, w_1231_, w_1707_);
and (w_0569_, new_in16[7], w_0579_);
not (w_0344_, w_0553_);
nand (w_0688_, new_in11[4], w_0781_);
nand (w_1203_, new_in13[5], new_in24[5]);
not (w_2093_, new_in10[8]);
xor (w_0247_, new_in5[0], new_in9[1]);
nand (w_1245_, w_0265_, w_0403_);
xor (w_0795_, new_in16[1], w_1839_);
and (w_1081_, w_1231_, w_0727_);
nand (w_1865_, new_in5[6], w_2205_);
nand (w_0409_, w_0742_, w_0696_);
xor (w_0140_, new_in16[1], w_0419_);
xor (w_2188_, new_in1[3], new_in8[2]);
xor (w_0107_, w_2109_, w_2149_);
xor (w_0711_, w_0150_, w_2167_);
or (w_1075_, w_2137_, w_0199_);
xor (w_1583_, w_0344_, w_2176_);
and (w_0186_, new_in20[0], w_0434_);
or (w_1829_, new_in1[1], w_1663_);
nand (w_2290_, new_in16[7], w_0863_);
nand (w_0610_, w_0923_, w_1082_);
xor (w_1549_, w_2195_, w_2257_);
nand (w_0146_, w_1231_, w_1643_);
or (w_1878_, w_0112_, w_2307_);
and (w_0872_, new_in5[6], w_0506_);
not (w_0441_, new_in13[2]);
xor (w_1493_, new_in3[3], w_1970_);
nand (w_1572_, w_1896_, w_0607_);
or (w_1260_, w_0958_, w_1865_);
nand (w_0386_, w_1253_, w_0957_);
nand (w_0907_, w_1011_, w_2309_);
nand (w_0547_, new_in17[1], new_in10[2]);
nand (w_1160_, w_0358_, w_0821_);
xor (w_0575_, w_0260_, w_1606_);
nand (w_0602_, new_in9[3], new_in15[3]);
nand (w_1677_, w_0581_, w_0348_);
or (w_0082_, w_2130_, w_1901_);
xor (w_1225_, w_0694_, w_1759_);
xor (w_1176_, new_in7[4], new_in15[4]);
nand (new_out13[4], w_1143_, w_1981_);
xor (w_2207_, new_in7[5], new_in15[5]);
nand (w_0125_, w_1151_, w_0500_);
xor (w_1618_, new_in1[1], new_in9[1]);
and (w_2273_, w_0719_, w_2164_);
xor (w_1748_, new_in4[4], w_1106_);
or (w_0154_, w_0539_, w_0935_);
xor (w_1576_, new_in22[2], w_0392_);
nand (w_1971_, w_0181_, w_1065_);
nand (w_0541_, w_2085_, w_2101_);
nand (w_1610_, w_1127_, w_0087_);
xor (w_0390_, new_in3[6], w_2019_);
nand (w_2058_, w_0707_, w_0734_);
xor (w_0343_, w_0165_, w_0444_);
nand (w_0652_, w_0244_, w_0826_);
nand (w_0682_, w_0250_, w_2097_);
xor (w_1563_, new_in23[0], new_in6[0]);
nand (w_0899_, w_1953_, w_1763_);
nand (w_1975_, w_1815_, w_2079_);
nand (w_1863_, w_1150_, w_1057_);
and (w_1575_, w_0508_, w_0294_);
and (w_1554_, w_0584_, w_1519_);
xor (w_1800_, new_in7[2], new_in15[2]);
or (w_0007_, w_1265_, w_2118_);
nand (w_0903_, w_0923_, w_1662_);
xor (w_1673_, w_1452_, w_0359_);
xor (w_1074_, w_0200_, w_2095_);
xor (w_0823_, w_1011_, w_0549_);
nor (w_1983_, w_0263_, w_0658_);
xor (w_1438_, w_0944_, w_0847_);
xor (w_0294_, w_0318_, w_0047_);
xor (w_1156_, new_in6[2], new_in18[2]);
and (w_1767_, w_1231_, w_0277_);
xor (w_2139_, new_in20[2], new_in11[2]);
or (w_0474_, w_2144_, w_1703_);
or (w_1105_, w_0789_, w_1674_);
nand (w_0317_, w_0168_, w_2316_);
or (w_0662_, w_0759_, w_0005_);
and (w_1344_, w_0263_, w_0720_);
or (w_1682_, w_0988_, w_1458_);
nand (w_1072_, w_1428_, w_0373_);
xor (w_1352_, new_in19[6], new_in17[6]);
nand (w_0057_, w_0725_, w_0167_);
xor (w_1363_, w_1853_, w_1599_);
nand (w_0578_, new_in16[3], w_0293_);
and (w_0995_, new_in18[0], new_in6[1]);
nand (w_1600_, w_1331_, w_1571_);
nand (w_1787_, w_0754_, w_2283_);
xor (w_0208_, w_0381_, w_2297_);
xor (w_1822_, w_0357_, w_1616_);
nand (w_1287_, w_0067_, w_0042_);
nand (w_1717_, new_in16[0], w_1343_);
xor (w_1533_, w_2007_, w_1126_);
nand (w_0073_, w_0730_, w_0904_);
xor (w_1030_, w_1365_, w_0314_);
or (w_2075_, w_0263_, w_0176_);
nand (w_1399_, w_0200_, w_2095_);
nand (w_0789_, new_in10[8], w_0263_);
xor (w_0581_, new_in9[0], new_in15[0]);
nand (w_0205_, w_0759_, w_0005_);
or (w_1266_, w_1538_, w_1585_);
nand (w_1667_, w_1835_, w_1285_);
nand (w_0416_, w_1234_, w_1788_);
and (w_1591_, w_1890_, w_1518_);
and (w_1685_, w_1423_, w_0575_);
nand (w_1488_, new_in16[3], w_1650_);
nand (new_out15[4], w_0028_, w_1241_);
and (w_0794_, w_0923_, w_0013_);
or (w_0454_, w_1427_, w_0245_);
xor (w_2271_, w_1670_, w_0471_);
xor (w_0284_, w_1596_, w_1268_);
or (w_1304_, w_1231_, w_0917_);
xor (w_1952_, w_0534_, w_1565_);
and (w_1515_, w_0630_, w_2017_);
nand (w_1296_, new_in12[1], new_in22[1]);
xor (w_0810_, new_in15[4], new_in9[4]);
nand (w_0902_, w_1717_, w_0140_);
or (w_0123_, new_in19[5], new_in17[5]);
xor (w_0848_, new_in7[5], new_in14[5]);
or (w_0234_, w_0091_, w_1140_);
or (w_1490_, w_1716_, w_1984_);
or (w_2103_, w_0263_, w_1416_);
or (w_0839_, w_0267_, w_1804_);
nand (w_1150_, w_0881_, w_1004_);
xor (w_1202_, w_0922_, w_1464_);
or (w_0959_, w_1231_, w_0792_);
xor (w_0749_, new_in20[1], new_in11[1]);
nand (w_1594_, new_in16[7], w_1598_);
xor (w_2057_, w_2235_, w_1022_);
and (w_0492_, w_2291_, w_2020_);
or (w_0858_, w_1315_, w_1107_);
xor (w_0053_, w_1619_, w_1256_);
or (w_0798_, w_1116_, w_2186_);
nand (w_1494_, w_1619_, w_1678_);
nand (w_2173_, w_1234_, w_0046_);
xor (w_0746_, w_0560_, w_0791_);
or (w_1669_, w_0091_, w_0893_);
xor (w_0445_, w_0121_, w_0626_);
nand (w_0819_, new_in20[4], w_1781_);
nand (w_0864_, new_in22[2], new_in14[1]);
or (w_2205_, w_0773_, w_1238_);
nand (w_1324_, w_0750_, w_1353_);
nand (new_out1[4], w_1421_, w_1163_);
nand (w_1570_, w_1967_, w_1360_);
nand (w_1037_, new_in10[8], w_0256_);
xor (w_0147_, new_in16[0], w_0244_);
and (w_2258_, w_0263_, w_2221_);
nand (w_0058_, w_0283_, w_0822_);
xor (w_1876_, w_0988_, w_1458_);
nand (w_0937_, w_2298_, w_0379_);
nand (w_2150_, w_1484_, w_0509_);
and (w_0055_, w_0263_, w_0898_);
and (new_out17[3], w_2094_, w_1303_);
and (w_0239_, w_0263_, w_0812_);
nand (w_0370_, w_1728_, w_1645_);
and (w_2238_, new_in10[8], w_0632_);
nand (w_1658_, w_1231_, w_1235_);
or (w_1736_, new_in8[0], w_1467_);
not (w_0006_, w_1250_);
nand (w_0645_, w_1968_, w_1430_);
xor (w_1729_, w_1191_, w_0976_);
nand (w_0866_, w_0972_, w_0908_);
and (w_1209_, new_in12[2], new_in15[0]);
nand (w_2113_, new_in16[2], w_1202_);
nand (w_0740_, w_0136_, w_0007_);
nand (w_0612_, new_in13[4], new_in24[4]);
xor (w_0982_, w_0114_, w_0287_);
and (new_out7[2], w_0552_, w_0157_);
nand (w_1526_, new_in5[6], w_0325_);
xor (w_2121_, new_in1[0], new_in9[0]);
xor (w_1980_, w_2085_, w_2101_);
nand (w_0528_, w_2093_, w_1054_);
nand (w_0309_, new_in19[2], new_in17[2]);
xor (w_1441_, new_in22[0], new_in21[0]);
and (w_2307_, w_1966_, w_1971_);
nand (w_0181_, w_0969_, w_0853_);
and (w_1331_, w_1231_, w_0923_);
or (w_1060_, w_2001_, w_2255_);
nand (w_1171_, w_0921_, w_1894_);
and (w_2131_, w_0923_, w_0820_);
xor (w_1107_, new_in22[5], w_0199_);
or (w_0577_, w_1214_, w_1801_);
or (w_1077_, w_0263_, w_1048_);
nand (w_2016_, w_1272_, w_1043_);
xor (w_0306_, w_1275_, w_1164_);
nand (w_0805_, w_1960_, w_0584_);
nand (w_1659_, w_0263_, w_1742_);
nand (w_1261_, w_1231_, w_1787_);
nand (w_2080_, new_in4[3], new_in2[3]);
xor (w_2208_, w_2067_, w_0828_);
and (w_0954_, w_0923_, w_1907_);
and (w_0696_, new_in5[6], w_1872_);
xor (w_0197_, new_in14[4], new_in22[5]);
nand (w_1419_, w_1843_, w_0163_);
xor (w_1279_, new_in24[5], new_in2[5]);
nand (w_1169_, w_1905_, w_0294_);
xor (w_1460_, w_1777_, w_1818_);
and (w_0669_, w_0951_, w_1293_);
nand (w_0508_, w_1571_, w_1314_);
xor (w_0663_, new_in14[4], new_in22[4]);
nand (w_2018_, w_0943_, w_0014_);
nand (w_0980_, new_in16[7], w_1868_);
nand (new_out14[1], w_1600_, w_0839_);
nand (w_0586_, w_0165_, w_0444_);
and (w_1099_, w_1231_, w_0391_);
or (w_1220_, w_1231_, w_0385_);
xor (w_1684_, new_in12[4], new_in15[2]);
xor (w_1624_, w_0482_, w_1748_);
xor (w_0784_, w_1491_, w_1424_);
xor (w_0653_, w_2070_, w_0845_);
nand (w_2094_, w_2093_, w_1760_);
nand (w_1178_, w_0534_, w_1565_);
nand (w_0157_, w_0004_, w_1655_);
or (w_0222_, w_1100_, w_1492_);
xor (w_1703_, new_in13[1], new_in1[1]);
nand (w_1535_, w_0121_, w_0626_);
nand (w_2089_, new_in5[2], new_in9[3]);
xor (w_0210_, new_in24[1], new_in2[1]);
nand (w_1227_, w_0205_, w_1632_);
and (w_0369_, new_in10[8], w_0231_);
and (w_1092_, new_in12[0], new_in19[0]);
or (w_0776_, w_0263_, w_2242_);
nand (new_out12[2], w_1142_, w_1323_);
nand (w_0279_, w_1231_, w_1660_);
xor (w_0036_, w_1537_, new_in12[4]);
xor (w_0826_, new_in21[0], new_in3[0]);
nand (w_1325_, w_0382_, w_0238_);
xor (w_0516_, new_in21[2], new_in3[2]);
and (w_1282_, new_in23[1], new_in12[1]);
nand (w_2046_, new_in19[3], new_in12[3]);
nand (w_1236_, new_in18[3], new_in6[4]);
nand (w_0712_, w_1462_, w_0088_);
nand (w_0420_, w_1372_, w_0443_);
xor (w_0633_, w_1415_, w_0669_);
xor (w_1851_, w_0514_, w_0081_);
nand (w_1836_, w_0129_, w_0350_);
xor (w_1407_, new_in16[4], w_1440_);
nand (w_1955_, new_in16[1], w_0887_);
nor (new_out12[3], w_1912_, w_0166_);
or (w_2212_, w_0263_, w_1946_);
and (w_1479_, w_2089_, w_0191_);
xor (w_1812_, w_0368_, w_1740_);
xor (w_1004_, new_in14[1], new_in21[1]);
xor (w_0287_, new_in17[1], new_in10[1]);
or (w_1730_, w_2145_, w_0981_);
nand (w_1394_, w_2117_, w_0802_);
nand (new_out5[1], w_1676_, w_1620_);
xor (w_1759_, w_0401_, w_0848_);
or (w_1968_, w_2124_, w_1273_);
not (w_2175_, w_1311_);
nand (w_0990_, new_in5[6], w_1429_);
nor (new_out1[3], w_1358_, w_2258_);
nand (w_1688_, new_in8[0], new_in5[6]);
nand (w_0716_, w_1838_, w_1755_);
xor (w_1120_, new_in14[1], new_in22[1]);
nand (w_0487_, w_2093_, w_0596_);
or (w_2021_, w_0422_, w_1563_);
nand (w_2279_, w_0998_, w_1410_);
and (new_out8[4], w_1454_, w_0930_);
xor (w_0583_, w_1875_, w_1383_);
not (w_0414_, w_0773_);
and (new_out17[0], w_1028_, w_0566_);
or (w_1076_, w_0567_, w_2281_);
xor (w_0471_, new_in4[1], new_in3[1]);
nand (w_0989_, w_1702_, w_1706_);
and (w_0326_, w_0913_, w_0342_);
or (w_1049_, w_1326_, w_0559_);
xor (w_0453_, w_0769_, w_1583_);
not (w_1537_, new_in23[4]);
nand (w_2191_, w_1139_, w_0259_);
xor (w_1435_, w_0943_, w_0151_);
xor (w_0705_, w_2284_, w_0460_);
and (w_0429_, w_0798_, w_2077_);
nand (w_1391_, w_0114_, w_0287_);
or (w_0108_, w_0680_, w_0672_);
nand (w_0707_, w_0075_, w_2185_);
nand (w_0405_, new_in4[1], w_0860_);
nand (w_1501_, w_1231_, w_0835_);
nand (w_1165_, w_1238_, w_2309_);
nand (w_1862_, new_in5[6], w_1161_);
xor (w_0726_, new_in20[1], w_1673_);
nand (w_1784_, w_1234_, w_1798_);
nand (w_1556_, w_0923_, w_1877_);
and (w_1683_, w_0263_, w_0682_);
nand (w_0277_, w_1322_, w_0593_);
or (w_0400_, w_1232_, w_1780_);
nand (new_out13[6], w_0461_, w_2082_);
xor (w_2176_, new_in1[5], new_in9[5]);
and (w_0136_, w_0263_, new_in5[6]);
nand (w_1109_, w_1297_, w_0555_);
or (w_0065_, w_0228_, w_0416_);
and (new_out9[2], w_0537_, w_1639_);
and (new_out17[4], w_1652_, w_2304_);
nand (w_1561_, w_2058_, w_0756_);
nand (w_1855_, w_0263_, w_0364_);
and (w_1654_, w_0923_, w_0469_);
xor (w_2306_, w_0609_, w_1357_);
and (w_0426_, new_in7[0], new_in8[1]);
and (w_0567_, new_in23[0], new_in6[0]);
xor (w_0489_, new_in1[0], new_in1[1]);
xor (w_1705_, new_in7[0], new_in8[1]);
xor (w_1527_, new_in11[6], new_in18[6]);
xor (w_1154_, w_0937_, w_0145_);
and (w_0668_, w_1785_, w_0484_);
xor (w_1719_, w_0036_, w_1284_);
or (w_2112_, new_in5[2], new_in9[3]);
and (w_1334_, w_1376_, w_1348_);
xor (w_0485_, w_0797_, w_1176_);
xor (w_1781_, w_0592_, w_0686_);
and (w_0144_, new_in20[0], w_2198_);
and (w_0085_, new_in16[7], w_1668_);
nand (w_0083_, w_1647_, new_in17[5]);
xor (w_1301_, new_in21[5], new_in20[6]);
nand (w_1495_, new_in7[2], new_in15[2]);
xor (w_0040_, new_in22[2], w_0871_);
or (w_1773_, w_0091_, w_0867_);
nand (w_2234_, w_0423_, w_1019_);
nand (w_1012_, w_1234_, w_1723_);
nand (w_2067_, w_0206_, w_0304_);
nor (w_1518_, new_in10[8], new_in5[6]);
or (w_0320_, w_1231_, w_2249_);
xor (w_1128_, new_in4[1], new_in2[1]);
and (w_0158_, new_in12[0], new_in22[0]);
and (w_1978_, w_1905_, w_0588_);
nand (w_0238_, w_0050_, w_0749_);
nand (w_1939_, new_in5[6], new_in7[0]);
nand (w_2182_, new_in22[4], new_in9[1]);
nand (w_1233_, w_1231_, w_0761_);
nor (w_2231_, w_0695_, new_in12[3]);
nand (new_out9[0], w_0472_, w_0064_);
xor (w_0042_, w_1613_, w_0625_);
nand (w_1032_, new_in1[1], new_in8[1]);
or (w_1413_, w_1231_, w_0581_);
xor (w_1795_, w_0384_, w_0849_);
nand (w_1252_, new_in7[3], new_in7[2]);
nand (w_1653_, w_0678_, w_1036_);
nand (w_1058_, w_1995_, w_1987_);
and (w_0809_, w_1000_, w_1944_);
xor (w_0791_, new_in17[1], new_in10[2]);
or (w_2286_, w_1791_, w_0051_);
nand (w_0072_, w_1231_, w_0303_);
nand (w_1053_, new_in5[6], w_0605_);
xor (w_2149_, new_in12[6], new_in15[4]);
nand (w_0974_, w_1753_, w_0137_);
nand (w_2264_, w_0864_, w_0693_);
xor (w_2198_, new_in10[0], new_in17[0]);
nand (w_1958_, w_2057_, w_2208_);
and (w_2254_, new_in5[6], w_1114_);
nand (w_0486_, new_in19[3], new_in6[2]);
and (w_2143_, w_1018_, w_1547_);
xor (w_2216_, w_0202_, w_1368_);
xor (w_1329_, new_in16[4], w_2147_);
and (w_0166_, w_1842_, w_2289_);
nand (w_1741_, w_1477_, w_0871_);
nand (w_0230_, w_1231_, w_0709_);
or (w_2069_, new_in18[2], new_in6[3]);
nand (w_0439_, w_1085_, w_0687_);
and (w_1213_, w_2093_, w_1060_);
xor (w_0790_, w_0459_, w_1110_);
xor (w_0699_, w_1318_, w_2015_);
nand (w_2233_, w_0992_, w_0532_);
and (new_out3[3], w_1754_, w_2268_);
nand (w_2136_, new_in7[3], new_in8[4]);
and (w_0706_, w_1905_, w_0718_);
xor (w_0188_, w_1419_, w_0481_);
not (w_0564_, w_1576_);
xor (w_1909_, w_1011_, w_2309_);
and (new_out7[3], w_2075_, w_0404_);
nand (w_2213_, new_in5[6], w_0603_);
nand (w_2125_, w_0129_, w_1188_);
and (w_1263_, new_in5[6], w_0130_);
and (w_1670_, new_in4[0], new_in3[0]);
nand (w_0148_, w_0788_, w_0606_);
nand (w_0500_, w_1290_, w_1066_);
xor (w_1013_, w_1834_, w_1527_);
or (w_0767_, w_2093_, w_0938_);
nand (w_0178_, w_1209_, w_2120_);
xor (w_0736_, new_in9[3], new_in15[3]);
nand (w_0424_, new_in1[0], w_0136_);
xor (w_1555_, w_0642_, w_1509_);
xor (w_0090_, new_in7[3], new_in7[2]);
and (w_1938_, w_1075_, w_0858_);
and (w_1957_, w_2011_, w_0910_);
nand (w_0312_, w_1427_, w_0290_);
nand (w_1999_, w_2093_, w_1459_);
nand (w_0727_, new_in10[0], w_1234_);
nand (w_1319_, new_in4[1], new_in2[1]);
or (w_0603_, new_in13[0], new_in1[0]);
nand (w_0945_, w_0188_, w_1604_);
nand (w_1691_, new_in5[6], w_2169_);
nand (w_0371_, new_in16[7], w_1747_);
nand (w_0531_, w_0507_, new_in17[1]);
nand (w_0536_, w_1330_, w_1599_);
xor (w_1031_, w_2084_, w_1812_);
nand (w_1676_, w_2200_, w_1764_);
nand (w_0468_, new_in18[1], new_in20[2]);
xor (w_0151_, w_0730_, w_0904_);
nand (w_1517_, w_2010_, w_2172_);
or (w_1041_, w_1038_, w_1881_);
xor (w_1145_, w_1113_, w_0396_);
xor (w_1354_, w_1995_, w_0319_);
xor (w_1899_, w_1637_, w_1492_);
xor (w_1064_, new_in20[2], w_0975_);
or (w_0248_, w_1231_, w_2051_);
nand (w_2268_, w_2093_, w_0764_);
nand (w_1609_, w_1991_, w_2050_);
nand (new_out16[4], w_0347_, w_2000_);
nand (w_1412_, w_0486_, w_0782_);
xor (w_2224_, w_0138_, w_0765_);
and (w_1126_, new_in23[5], new_in12[5]);
and (w_1846_, w_1441_, w_0546_);
nand (w_2128_, w_0932_, w_0902_);
nand (w_0833_, w_1905_, w_2141_);
nand (w_0987_, new_in20[1], w_1673_);
or (w_0496_, w_0929_, w_0906_);
xor (w_0385_, w_0678_, w_1036_);
and (w_1351_, new_in16[7], w_1996_);
nand (new_out3[0], w_1999_, w_1734_);
nand (w_0921_, new_in14[3], new_in22[4]);
and (new_out6[0], w_2087_, w_1335_);
and (w_1525_, w_0286_, w_1710_);
xor (w_1461_, w_1253_, w_0957_);
nand (new_out4[3], w_0948_, w_0279_);
nor (w_0278_, w_1567_, w_0218_);
and (w_1582_, new_in14[0], new_in22[1]);
nand (w_0138_, w_1921_, w_1636_);
or (w_0334_, w_1677_, w_0470_);
nor (new_out11[1], w_1983_, w_0399_);
xor (w_1961_, new_in9[1], new_in15[1]);
xor (w_0033_, w_1202_, w_2259_);
xor (w_2190_, w_1689_, w_0210_);
and (w_1234_, new_in10[8], w_0263_);
nand (w_0888_, w_1574_, w_2197_);
xor (w_1521_, new_in19[2], new_in12[2]);
xor (w_1700_, new_in13[2], new_in24[2]);
xor (w_2185_, w_1962_, w_1534_);
and (w_0237_, new_in10[8], w_0841_);
and (w_1530_, w_1687_, w_2116_);
and (w_0912_, w_2055_, w_2036_);
nand (w_1833_, w_1738_, w_1618_);
xor (w_1910_, w_1728_, w_1645_);
nand (new_out2[1], w_0834_, w_2150_);
xor (w_1048_, new_in9[0], w_0247_);
xor (w_1177_, w_0655_, w_0575_);
nand (w_1364_, w_2282_, w_0262_);
nand (w_2298_, new_in1[4], new_in8[4]);
xor (w_0176_, w_0132_, w_0704_);
xor (w_0599_, w_1527_, w_0492_);
xor (w_0005_, w_2171_, w_1515_);
nand (w_0190_, w_1500_, w_1906_);
or (w_1118_, w_0186_, w_0726_);
or (w_0762_, w_1405_, w_1576_);
xor (w_1050_, w_1442_, w_0264_);
xor (w_1123_, new_in14[5], new_in21[5]);
nand (w_0043_, w_1880_, w_0897_);
nand (w_2110_, w_1231_, w_0753_);
or (w_0463_, w_0283_, w_0833_);
xor (w_0561_, new_in19[0], new_in19[1]);
nand (w_1442_, w_0634_, w_2162_);
xor (w_0781_, w_0870_, w_1672_);
or (w_2030_, w_1507_, w_0209_);
xor (w_0490_, w_2026_, w_1585_);
and (w_2007_, w_0609_, w_1357_);
or (w_1223_, w_0263_, w_1557_);
xor (w_2138_, w_0775_, w_2016_);
and (w_1211_, w_1133_, w_2266_);
nand (w_0654_, w_1095_, w_1153_);
and (w_1916_, w_1972_, w_1003_);
or (w_0862_, w_1231_, w_2121_);
nand (w_1849_, w_1373_, w_1712_);
and (w_1644_, w_1287_, w_1072_);
xor (w_1881_, w_0637_, w_2207_);
nand (w_1859_, w_2159_, w_0570_);
or (w_1278_, w_1769_, w_0020_);
xor (w_1948_, w_1991_, w_2050_);
and (w_0940_, new_in16[7], w_0836_);
xor (w_0685_, w_0125_, w_1593_);
nand (w_1020_, w_1419_, w_0481_);
nand (w_2119_, new_in19[1], new_in17[1]);
not (w_1647_, new_in19[5]);
nand (w_1724_, w_0144_, w_1891_);
nand (w_0459_, new_in23[2], new_in12[2]);
xor (w_2041_, new_in21[1], new_in3[1]);
and (w_1528_, w_0632_, w_1210_);
nand (w_0587_, new_in16[7], w_0939_);
or (w_2053_, new_in19[3], w_1401_);
xor (w_1369_, w_2099_, w_2040_);
nand (w_0527_, w_0553_, w_2176_);
xor (w_1951_, w_0911_, w_0647_);
nand (w_1746_, w_1083_, w_1829_);
nand (w_0730_, w_1915_, w_0089_);
nand (w_1885_, w_2214_, w_2202_);
nand (w_0008_, new_in1[2], new_in8[2]);
and (w_0228_, w_1820_, w_2038_);
nand (w_0638_, w_1304_, w_0805_);
nor (w_0883_, w_1769_, w_0020_);
xor (w_2301_, w_1993_, w_0777_);
xor (w_1267_, w_0168_, w_2316_);
and (w_2135_, w_0370_, w_0299_);
nand (w_0753_, w_1866_, w_0027_);
xor (w_1385_, new_in16[5], w_0199_);
xor (w_1945_, w_2102_, w_0242_);
xor (w_1623_, w_1790_, w_1864_);
nand (w_0406_, w_1614_, w_1914_);
and (w_1695_, new_in5[2], w_0601_);
nand (w_0292_, new_in8[1], w_0994_);
xor (w_1559_, w_0892_, w_1590_);
xor (w_0249_, w_1530_, w_0589_);
or (w_1395_, w_1817_, w_0783_);
nand (w_0174_, w_0574_, w_1584_);
nand (w_0351_, w_0056_, w_1761_);
and (w_1678_, new_in5[6], w_1041_);
and (w_2232_, w_1545_, w_0488_);
nand (w_1708_, new_in11[3], w_2181_);
xor (w_2157_, new_in1[0], w_2056_);
nand (w_1111_, w_1453_, w_1961_);
nand (w_1715_, new_in21[4], new_in3[4]);
nand (w_1707_, new_in19[0], w_1234_);
nand (w_0472_, w_1413_, w_0055_);
xor (w_0361_, new_in20[0], w_0434_);
nand (w_1045_, w_1251_, w_0369_);
or (w_0985_, w_0263_, w_1624_);
xor (w_1884_, new_in18[4], new_in6[5]);
xor (w_1482_, w_2166_, w_1014_);
xor (w_1159_, w_1100_, w_1492_);
nand (w_1832_, new_in19[4], new_in17[4]);
and (w_2230_, new_in5[6], w_0388_);
nand (w_1232_, w_2093_, new_in16[7]);
nand (w_0120_, w_0497_, w_1162_);
nand (w_2066_, new_in1[3], new_in13[3]);
or (w_1574_, w_2093_, w_0561_);
and (w_0110_, w_2245_, w_1731_);
and (w_1651_, w_2178_, w_1827_);
nand (w_1087_, w_1503_, w_0258_);
nand (w_2055_, new_in22[1], w_0887_);
nand (w_1699_, new_in7[1], new_in8[2]);
not (w_2237_, w_0906_);
xor (w_2090_, new_in21[4], new_in20[5]);
nand (w_0799_, new_in16[7], w_2252_);
xor (w_1082_, w_1278_, w_1141_);
nand (w_0996_, new_in4[4], new_in2[4]);
nand (w_0905_, w_1231_, w_1711_);
nand (new_out12[1], w_0834_, w_1932_);
and (w_1740_, w_0949_, w_1936_);
and (w_1427_, new_in22[0], new_in16[0]);
and (w_2221_, w_1185_, w_1149_);
nand (w_1468_, w_2260_, w_1686_);
or (w_0265_, w_2145_, w_0544_);
xor (w_2252_, w_1447_, w_0656_);
nand (w_1008_, w_1543_, w_0276_);
and (w_1281_, w_1905_, w_0417_);
nand (w_1138_, w_1231_, w_2238_);
xor (w_0934_, w_0758_, w_1173_);
nand (w_1898_, w_1180_, w_0999_);
nand (w_0874_, new_in20[3], new_in11[3]);
or (w_0629_, w_0324_, w_0479_);
xor (w_0860_, w_0844_, w_2155_);
xor (w_1911_, w_1634_, w_0550_);
xor (w_2095_, w_0800_, w_2321_);
nand (w_0757_, new_in7[4], new_in15[4]);
nand (w_0347_, w_1023_, w_1277_);
xor (w_1210_, w_1325_, w_2139_);
nand (w_0747_, w_0559_, w_1019_);
nand (w_0524_, new_in9[1], new_in15[1]);
nand (w_0340_, w_1347_, w_1356_);
xor (w_1472_, new_in7[3], new_in8[4]);
xor (w_2050_, new_in20[3], new_in11[3]);
nand (w_1792_, w_0573_, w_1771_);
not (w_1398_, new_in13[1]);
or (w_0296_, w_0263_, w_1267_);
xor (w_0086_, w_1750_, w_1337_);
xor (w_1390_, w_1964_, w_0895_);
and (w_0135_, w_0263_, w_1504_);
and (w_0594_, w_2097_, w_1511_);
xor (w_1280_, new_in22[2], new_in14[2]);
xor (w_2034_, w_1519_, w_2157_);
nand (w_0963_, new_in5[6], w_1422_);
nand (w_1696_, new_in1[3], new_in8[3]);
nand (w_0563_, w_0771_, w_1940_);
nand (w_0731_, w_0186_, w_0726_);
nand (w_0064_, new_in16[7], w_0501_);
nand (w_1434_, new_in5[6], w_1154_);
nand (w_0715_, w_1204_, w_0721_);
or (w_1429_, w_0958_, w_2048_);
nand (w_1713_, new_in23[2], new_in6[2]);
and (w_0088_, new_in5[6], w_0474_);
xor (w_2181_, w_0407_, w_0225_);
xor (w_0204_, w_1063_, w_1206_);
or (w_1079_, w_1582_, w_1692_);
nand (w_0744_, w_1956_, w_2192_);
xor (w_2040_, w_0717_, w_1800_);
nand (w_2280_, new_in19[4], new_in6[3]);
xor (w_0015_, new_in13[4], new_in1[4]);
xor (w_0703_, new_in17[4], new_in10[5]);
xor (w_0348_, new_in13[0], new_in24[0]);
nand (w_0593_, w_0652_, w_2131_);
nand (w_1127_, w_0923_, w_1435_);
nand (w_0000_, w_0909_, w_1860_);
and (w_0616_, new_in12[0], new_in23[0]);
nand (new_out13[3], w_1658_, w_2133_);
xor (w_1359_, new_in5[1], new_in9[2]);
xor (w_1119_, new_in1[2], new_in8[1]);
nand (w_1888_, new_in16[1], w_1839_);
or (w_1023_, w_0263_, w_1144_);
and (w_1423_, w_0944_, w_1363_);
nand (w_1292_, w_0410_, w_1554_);
xor (w_0734_, w_1900_, w_1274_);
xor (w_1723_, w_1628_, w_1816_);
not (w_1231_, new_in5[6]);
nand (w_0565_, w_2274_, w_2188_);
nand (w_0924_, w_1231_, w_0814_);
and (new_out6[2], w_0840_, w_1245_);
nand (w_0493_, w_0188_, w_1951_);
and (w_0919_, w_1388_, w_1821_);
nand (w_0875_, w_0263_, w_0888_);
xor (w_1940_, new_in1[3], new_in13[3]);
or (w_1305_, w_1231_, w_0955_);
nand (w_1098_, new_in10[8], w_1922_);
xor (w_1589_, new_in6[3], new_in18[3]);
and (new_out15[2], w_0799_, w_1371_);
and (w_0570_, w_0923_, w_2174_);
nand (w_0686_, w_1196_, w_1061_);
and (w_1538_, w_1198_, w_1183_);
xor (w_0773_, w_1453_, w_1961_);
nand (w_1474_, new_in19[3], w_1401_);
nand (w_1564_, new_in20[2], new_in11[2]);
and (w_0584_, new_in16[7], w_1231_);
nand (w_1194_, new_in18[4], new_in11[4]);
xor (w_1317_, w_0633_, w_0355_);
and (w_1627_, w_0879_, w_1134_);
nand (w_2177_, w_0995_, w_1690_);
and (w_1580_, w_1830_, w_0454_);
nand (w_2123_, w_0263_, w_1698_);
nand (w_0193_, w_1318_, w_2015_);
or (w_0175_, w_1964_, w_0895_);
xor (w_1144_, w_2206_, w_2170_);
nand (w_0102_, w_1558_, w_1024_);
xor (w_1765_, new_in20[4], new_in11[4]);
or (w_1866_, w_2093_, w_2323_);
nand (w_1093_, w_1053_, w_0582_);
or (w_1830_, w_0789_, w_2198_);
xor (w_0556_, w_1901_, w_1384_);
xor (w_2051_, new_in22[0], w_0861_);
nand (w_2160_, w_1836_, w_0104_);
nand (w_0308_, w_1716_, w_1984_);
and (w_1982_, w_0451_, w_1994_);
and (w_1090_, new_in16[7], w_0615_);
nand (w_1941_, w_0266_, w_1281_);
xor (w_0246_, new_in12[0], new_in23[0]);
nand (w_0738_, w_1495_, w_0039_);
nand (new_out18[6], w_0116_, w_1217_);
xor (w_1508_, new_in22[2], w_0733_);
nand (w_2004_, w_0748_, w_1521_);
and (w_1137_, new_in10[8], w_1377_);
xor (w_0765_, w_1647_, new_in12[5]);
xor (w_1807_, new_in4[4], new_in3[4]);
nand (w_1687_, new_in9[5], new_in15[5]);
xor (w_0397_, w_1701_, w_0698_);
or (w_1919_, w_0263_, w_0970_);
nand (w_2153_, w_0083_, w_0993_);
nand (w_0382_, new_in20[1], new_in11[1]);
xor (w_1606_, new_in1[4], new_in9[4]);
and (w_0118_, w_1258_, w_2236_);
or (w_1046_, w_1357_, w_0362_);
xor (w_0423_, w_1008_, w_0201_);
nand (w_0702_, w_0408_, w_1808_);
xor (w_0020_, w_0158_, w_1417_);
and (w_1791_, w_0182_, w_1266_);
nand (w_1959_, w_2093_, w_1885_);
and (w_0701_, w_2209_, w_1099_);
or (w_0615_, w_1582_, w_0571_);
nor (w_1328_, w_0263_, w_0183_);
and (w_1906_, w_0263_, w_0675_);
nand (w_0596_, w_1305_, w_1292_);
xor (w_1789_, w_0431_, w_1588_);
nand (w_1235_, w_0857_, w_1803_);
nand (w_2043_, new_in5[6], w_0660_);
nand (w_2324_, w_1447_, w_0656_);
and (w_0114_, new_in10[0], new_in17[0]);
nand (w_1601_, w_0263_, w_1045_);
xor (w_0589_, new_in15[6], new_in9[6]);
and (w_1346_, w_0760_, w_0476_);
nand (w_0111_, w_0057_, w_1904_);
nand (w_0879_, new_in19[5], new_in6[4]);
nand (w_0323_, new_in7[3], new_in15[3]);
nand (w_1214_, w_1858_, w_0522_);
nand (w_0538_, w_1152_, w_0736_);
xor (w_1963_, new_in21[1], w_2001_);
nand (w_0023_, new_in18[3], new_in11[3]);
or (w_0739_, w_0789_, w_0876_);
nand (new_out4[4], w_0127_, w_0813_);
nand (w_1776_, w_1466_, w_0643_);
nand (new_out1[5], w_1379_, w_2134_);
nand (w_1635_, w_0044_, w_1855_);
nand (w_0211_, w_1378_, new_in17[2]);
xor (w_1588_, new_in18[4], new_in11[4]);
and (w_1874_, w_0991_, w_0446_);
nand (w_2033_, w_1905_, w_1869_);
xor (w_2244_, w_2232_, w_1135_);
nand (w_1136_, new_in16[7], w_1350_);
and (w_1453_, new_in9[0], new_in15[0]);
nand (w_0161_, w_0374_, w_2008_);
nand (w_2140_, w_2121_, w_0751_);
xor (w_2052_, new_in21[5], w_2078_);
nand (w_0315_, w_2012_, w_1062_);
xor (w_1404_, w_2057_, w_0648_);
xor (w_1770_, w_0096_, w_0067_);
and (w_0657_, w_1905_, w_1986_);
xor (w_0223_, w_1525_, w_2052_);
and (w_0591_, w_0263_, w_1448_);
nand (w_0949_, w_0800_, w_2057_);
and (w_0225_, w_1230_, w_2069_);
nand (w_1406_, new_in5[6], w_2163_);
and (w_1524_, new_in16[7], w_2003_);
and (new_out2[2], w_1142_, w_0928_);
or (w_1666_, w_2058_, w_0316_);
nand (w_0387_, w_0844_, w_2155_);
nand (w_0877_, new_in17[2], new_in10[2]);
nand (w_1573_, w_0227_, w_2045_);
xor (w_0268_, w_2282_, w_0262_);
xor (w_1743_, w_0079_, w_1407_);
xor (w_2027_, w_0884_, w_1029_);
nand (w_1091_, w_0228_, w_0150_);
nand (w_0333_, w_1243_, w_2004_);
nand (w_1714_, w_1894_, w_0010_);
nand (w_1987_, w_0778_, w_2119_);
or (w_0914_, w_0336_, w_1661_);
xor (w_1840_, w_0881_, w_0208_);
nor (new_out18[2], w_1328_, w_1333_);
nand (w_1372_, w_0568_, w_1068_);
nand (w_1504_, new_in5[6], w_1177_);
xor (w_0470_, w_0414_, w_0208_);
nand (w_2162_, w_1370_, w_1359_);
nand (w_0017_, new_in24[2], new_in2[2]);
nand (w_1481_, new_in10[8], w_1084_);
xor (w_1078_, w_2154_, w_1940_);
xor (w_1946_, w_1578_, w_1017_);
nand (w_0778_, w_1901_, w_1384_);
nand (w_2247_, w_1665_, w_0810_);
or (w_1907_, w_1512_, w_1965_);
nand (new_out6[4], w_1216_, w_1825_);
nand (w_2000_, new_in10[8], w_1948_);
xor (w_2179_, w_0965_, w_2090_);
and (w_1100_, w_2099_, w_2040_);
and (w_0977_, w_0263_, w_0177_);
or (w_0388_, w_1396_, w_0153_);
or (w_0011_, w_1828_, w_0012_);
nand (w_1571_, w_0802_, w_1076_);
nand (w_0365_, w_1234_, w_1822_);
or (w_1303_, w_2093_, w_0685_);
nand (w_0427_, w_0800_, w_2321_);
and (w_0679_, w_0211_, w_1121_);
and (w_1405_, w_1296_, w_1386_);
xor (w_0670_, w_2147_, w_0284_);
nand (w_1018_, new_in21[5], new_in3[5]);
nand (w_1921_, new_in19[4], new_in12[4]);
xor (w_1114_, new_in13[0], new_in5[0]);
and (new_out4[0], w_2246_, w_2083_);
nand (w_0671_, w_0120_, w_1288_);
xor (w_0735_, new_in20[0], new_in11[0]);
nand (w_2084_, w_0202_, w_0321_);
and (new_out18[0], w_0666_, w_0043_);
nand (w_0350_, w_1958_, w_1188_);
xor (w_0540_, new_in1[4], new_in8[3]);
nand (w_2287_, new_in22[4], w_2161_);
or (w_0618_, w_1231_, w_1990_);
and (w_1485_, w_2288_, w_1125_);
xor (w_1476_, w_1528_, w_1948_);
nand (w_2151_, w_1426_, w_1295_);
nand (w_1471_, w_1234_, w_0846_);
or (w_1668_, w_2264_, w_1621_);
nand (new_out3[4], w_0528_, w_1481_);
nand (w_0286_, new_in21[4], w_2303_);
xor (w_0012_, new_in12[1], w_0376_);
nand (w_1698_, w_1169_, w_2160_);
nand (w_2236_, w_2263_, w_0855_);
not (w_0600_, w_2010_);
nand (w_1375_, w_2166_, w_0623_);
xor (w_0024_, w_0110_, w_0933_);
nand (w_0475_, w_0398_, w_0119_);
nand (w_0328_, w_0423_, w_1249_);
nand (w_1540_, new_in16[7], new_in9[0]);
and (w_0741_, new_in7[2], new_in7[1]);
and (w_2145_, w_1522_, w_1310_);
nand (w_0172_, w_0230_, w_1526_);
nand (w_0574_, w_0031_, w_0308_);
xor (w_0664_, w_1478_, w_1743_);
xor (w_0893_, w_0115_, w_1751_);
xor (w_2146_, w_0715_, w_1472_);
nand (w_2211_, w_2292_, w_1349_);
xor (w_0155_, w_1307_, w_0679_);
nor (w_0950_, w_1470_, w_0151_);
or (w_0666_, w_0263_, w_1802_);
or (w_1149_, w_1231_, w_0311_);
xor (w_0887_, new_in23[1], w_0556_);
or (w_0604_, w_0263_, w_0851_);
nand (w_1858_, new_in14[2], new_in22[3]);
and (w_0649_, w_0115_, w_1751_);
or (w_0993_, w_1433_, w_1515_);
xor (w_1167_, new_in22[6], new_in9[3]);
xor (w_2323_, w_2314_, w_1963_);
nand (w_0745_, w_0694_, w_1759_);
or (w_1183_, w_0912_, w_1508_);
or (w_0691_, w_0144_, w_0035_);
or (w_2065_, w_1414_, w_2321_);
or (w_2283_, w_0263_, w_1497_);
xor (w_0785_, w_0995_, w_1690_);
nor (w_1513_, w_1231_, w_1316_);
nand (w_1181_, w_0650_, w_1239_);
nand (w_1071_, w_1696_, w_1181_);
xor (w_0512_, new_in24[4], new_in2[4]);
and (w_1339_, w_0263_, w_0942_);
nand (w_2005_, w_1294_, w_1244_);
nand (w_0200_, w_2037_, w_0317_);
nand (w_0281_, new_in12[5], new_in15[3]);
nand (w_1061_, w_0150_, w_2167_);
nand (w_2285_, new_in22[2], new_in16[2]);
nand (w_2178_, w_1340_, w_0954_);
xor (w_0016_, w_0340_, w_0194_);
nand (w_0241_, w_0700_, w_1645_);
and (w_0502_, w_0263_, w_2218_);
nand (w_0885_, w_2179_, w_1123_);
nand (new_out10[1], w_1115_, w_1908_);
xor (w_1798_, w_0931_, w_0703_);
nand (w_0998_, w_1425_, w_1896_);
nand (w_0523_, w_0881_, w_0208_);
nand (w_0031_, new_in20[3], w_0711_);
nand (w_2203_, new_in16[7], w_1441_);
nand (w_2255_, new_in16[7], w_1231_);
nand (w_2023_, w_0333_, w_0289_);
xor (w_1645_, w_0074_, w_1684_);
xor (w_1848_, w_1928_, w_1156_);
nand (w_1133_, new_in22[1], w_0376_);
nand (w_0624_, new_in5[6], w_1159_);
xor (w_0143_, new_in18[0], new_in6[1]);
nand (w_0233_, w_0911_, w_0647_);
xor (w_1157_, w_1732_, w_0829_);
and (w_1917_, w_0288_, w_2276_);
nand (w_0100_, w_0203_, w_1080_);
xor (w_1970_, w_1667_, w_0059_);
nand (w_0404_, w_1709_, w_1683_);
nand (w_1129_, new_in10[8], w_1848_);
and (w_1904_, new_in5[6], w_1224_);
xor (w_0466_, new_in13[5], new_in5[5]);
nand (new_out4[1], w_2110_, w_0409_);
and (w_1567_, new_in1[0], new_in1[1]);
nand (w_2049_, w_0965_, w_2090_);
nand (w_2199_, w_1905_, w_1851_);
xor (w_1337_, w_0741_, w_0090_);
and (w_1172_, w_0263_, w_0862_);
xor (w_0933_, w_0025_, w_0093_);
nand (w_1996_, w_1033_, w_1317_);
and (w_1229_, w_1148_, w_0878_);
nand (w_2012_, w_0920_, w_2032_);
and (w_1274_, w_0578_, w_0986_);
or (w_0588_, w_0616_, w_1282_);
nand (w_0562_, w_1446_, new_in7[4]);
xor (w_0259_, new_in18[2], new_in20[3]);
xor (w_0700_, new_in7[4], new_in14[4]);
nand (w_2024_, w_0614_, w_1854_);
nand (w_1190_, w_1234_, w_1845_);
or (w_1763_, w_2114_, w_0740_);
or (w_2158_, w_2093_, w_0359_);
xor (w_0221_, new_in17[3], new_in10[4]);
and (w_0723_, w_2064_, w_1020_);
nand (w_1811_, w_2093_, w_0172_);
nand (w_1896_, w_1817_, w_0783_);
nand (w_0947_, w_1332_, w_1724_);
xor (w_1690_, new_in18[1], new_in6[2]);
xor (w_1222_, new_in17[2], new_in10[3]);
xor (w_0105_, w_1930_, w_0235_);
and (w_2079_, w_1905_, w_0393_);
and (w_1927_, new_in8[0], new_in1[0]);
or (w_2091_, w_2198_, w_0287_);
nand (w_1389_, w_0773_, w_0208_);
xor (w_1492_, w_0738_, w_1697_);
nand (w_0078_, w_1190_, w_1531_);
xor (w_1854_, new_in11[4], w_0781_);
xor (w_2299_, w_0222_, w_0485_);
and (w_1808_, w_0263_, w_2187_);
xor (w_1175_, w_0030_, w_0491_);
xor (w_1164_, new_in24[6], new_in2[6]);
or (w_1646_, w_0735_, w_0422_);
nand (w_0231_, w_1627_, w_1300_);
or (w_0675_, w_2144_, w_2213_);
nand (w_0965_, w_0430_, w_0732_);
and (new_out8[2], w_0296_, w_1783_);
nand (w_0693_, w_1582_, w_0571_);
nand (w_1009_, w_0715_, w_1472_);
nand (w_2009_, new_in10[8], w_1539_);
xor (w_0183_, w_1863_, w_0823_);
nand (w_1914_, w_0381_, w_2297_);
xor (w_0041_, w_0439_, w_2215_);
xor (w_1239_, new_in1[3], new_in8[3]);
and (w_0421_, new_in10[8], w_1118_);
and (w_0264_, w_2089_, w_2112_);
xor (w_1796_, new_in7[6], new_in15[6]);
or (w_1892_, w_1231_, w_1806_);
nor (w_1630_, w_2168_, new_in17[3]);
xor (w_0884_, w_0390_, w_0723_);
not (w_1378_, new_in19[2]);
or (w_2003_, w_0147_, w_0494_);
nand (w_1330_, w_2220_, w_0152_);
or (w_0192_, w_0581_, w_0348_);
and (new_out1[0], w_0190_, w_2203_);
or (w_1349_, w_1231_, w_1770_);
nand (w_1817_, w_0405_, w_0997_);
xor (w_0850_, w_2048_, w_2208_);
nand (w_0598_, w_0111_, w_1949_);
or (w_0579_, w_1334_, w_0095_);
and (w_1511_, new_in13[0], new_in13[1]);
nand (w_1241_, new_in16[7], w_1552_);
nand (w_1421_, w_0263_, w_2310_);
nand (w_2267_, w_2035_, w_0330_);
nand (w_2266_, w_1925_, w_0070_);
nand (w_0035_, w_1905_, w_1929_);
xor (w_1542_, w_1355_, w_1805_);
and (w_0756_, new_in16[7], w_1969_);
nand (w_0395_, w_2145_, w_0981_);
and (w_1925_, new_in22[0], w_0861_);
xor (w_1368_, w_0825_, w_1498_);
or (w_2246_, w_1231_, w_1381_);
xor (w_0822_, new_in18[1], new_in20[2]);
nand (w_1257_, w_0520_, w_0516_);
or (w_1568_, w_0441_, w_0548_);
nand (w_1894_, w_1214_, w_1801_);
nand (w_0942_, w_0058_, w_1298_);
nand (w_1152_, w_1733_, w_2151_);
xor (w_2086_, new_in3[1], w_0811_);
nand (w_2159_, w_0713_, w_0670_);
xor (w_0251_, w_2012_, w_0934_);
nand (w_2193_, new_in19[1], new_in12[1]);
nand (w_0094_, w_1170_, w_0536_);
xor (w_0542_, new_in6[1], new_in18[1]);
or (w_0972_, w_1326_, w_0990_);
nand (w_1068_, w_0318_, w_0047_);
xor (w_1065_, new_in5[5], w_0708_);
or (w_0820_, w_0244_, w_0826_);
nand (w_2002_, w_0263_, w_2180_);
xor (w_1777_, new_in7[0], new_in15[0]);
or (w_1985_, w_2324_, w_1050_);
and (w_0052_, w_0796_, w_1546_);
nand (w_0936_, w_0437_, w_1178_);
nand (new_out10[4], w_0195_, w_0905_);
nand (w_1110_, w_0616_, w_1282_);
or (w_0832_, w_1578_, w_1017_);
nand (w_1856_, w_1231_, w_1841_);
nand (w_0650_, w_0008_, w_1653_);
xor (w_0311_, w_2249_, w_1078_);
nand (w_1016_, w_0112_, w_2307_);
nand (w_0720_, w_1905_, w_1533_);
xor (w_1439_, w_1982_, w_1611_);
and (w_0342_, w_1231_, w_1551_);
and (w_1085_, w_0049_, w_2146_);
nand (new_out10[2], w_1261_, w_0831_);
nand (w_0482_, w_1444_, w_2279_);
nand (w_0001_, new_in15[4], new_in9[4]);
xor (w_1844_, new_in21[6], new_in3[6]);
nand (w_1709_, w_1474_, w_2028_);
xor (w_1579_, w_2071_, w_2240_);
and (w_1353_, w_0263_, w_2021_);
xor (w_2305_, w_0049_, w_2146_);
nand (w_1403_, w_1905_, w_1207_);
nand (w_1462_, w_2144_, w_1703_);
xor (w_0915_, w_0181_, w_1065_);
nand (w_0030_, w_0817_, w_2275_);
xor (w_1739_, w_1201_, w_0249_);
not (w_1446_, new_in7[3]);
nand (w_0807_, w_1058_, w_0309_);
and (w_1779_, w_1905_, w_0467_);
nand (w_0550_, w_0441_, new_in13[3]);
nand (w_1734_, new_in10[8], w_0246_);
nand (w_1216_, w_1231_, w_1345_);
nand (w_1146_, w_0267_, w_1208_);
and (w_0988_, w_1741_, w_0842_);
nand (w_1566_, w_0523_, w_0354_);
or (w_1861_, w_0079_, w_1407_);
nand (w_1264_, w_0426_, w_2315_);
nand (w_0366_, w_0892_, w_1271_);
xor (w_1424_, w_1679_, w_0226_);
and (w_1893_, w_1941_, w_0077_);
nand (w_1094_, w_1613_, w_0625_);
nor (new_out5[5], w_1992_, w_0701_);
xor (w_0684_, new_in4[2], new_in3[2]);
xor (w_0606_, w_1238_, w_2309_);
and (w_0050_, new_in20[0], new_in11[0]);
nand (w_1466_, new_in19[2], new_in6[1]);
xor (w_0383_, new_in22[6], w_1308_);
xor (w_1457_, new_in18[3], new_in11[3]);
and (w_1401_, new_in19[2], w_0865_);
xor (w_1641_, w_2029_, w_0946_);
nand (w_1681_, w_1828_, w_0012_);
nand (new_out15[3], w_1025_, w_0702_);
nand (w_1083_, new_in1[0], w_0218_);
nand (w_0285_, new_in10[8], w_0735_);
and (w_0526_, w_0310_, w_0683_);
xor (w_0925_, new_in23[6], new_in6[6]);
xor (w_0845_, new_in18[4], new_in20[5]);
nand (w_1285_, w_2195_, w_2257_);
nand (w_1039_, new_in1[1], new_in9[1]);
xor (w_0824_, new_in1[1], new_in8[1]);
nand (w_1617_, new_in5[1], w_1487_);
xor (w_1522_, w_1427_, w_0290_);
nand (w_1028_, w_2093_, w_0638_);
nand (w_0495_, w_0096_, w_0113_);
nand (w_0156_, w_1566_, w_1909_);
nand (w_0109_, w_0691_, w_1172_);
and (w_1197_, new_in16[7], w_0692_);
xor (w_1005_, w_1242_, w_1807_);
xor (w_1069_, w_1189_, w_1597_);
or (w_0393_, w_0947_, w_1064_);
nand (w_2189_, w_0023_, w_2217_);
nand (w_1199_, w_1900_, w_0986_);
nand (w_0952_, w_0739_, w_1079_);
and (w_1333_, w_1431_, w_0591_);
xor (w_1104_, w_0395_, w_0511_);
nand (w_2322_, w_2147_, w_0284_);
or (w_0425_, w_2121_, w_0751_);
xor (w_1657_, new_in4[6], new_in2[6]);
nand (w_2167_, w_0877_, w_1675_);
nand (w_0021_, w_1556_, w_0029_);
xor (w_2320_, w_1047_, w_2301_);
xor (w_2319_, w_0936_, w_1974_);
nand (w_1170_, new_in1[3], new_in9[3]);
xor (w_0580_, new_in5[3], new_in9[4]);
nand (w_2156_, new_in9[0], new_in22[3]);
xor (w_0891_, w_0594_, w_0766_);
xor (w_1067_, w_1071_, w_0269_);
xor (w_1672_, new_in18[3], new_in6[4]);
nand (w_1890_, new_in16[7], w_1950_);
nand (w_2014_, w_1483_, w_2111_);
nand (w_0951_, new_in11[5], w_0525_);
nand (w_1686_, new_in10[8], w_1059_);
and (w_0667_, w_1083_, w_1086_);
nand (w_1614_, new_in13[1], new_in24[1]);
xor (w_1611_, new_in17[6], new_in10[6]);
xor (w_0957_, w_1520_, w_1735_);
or (w_0415_, w_2093_, w_1595_);
nand (w_0422_, new_in10[8], w_1231_);
or (w_0213_, w_1814_, w_2042_);
xor (w_2115_, w_2065_, w_1645_);
xor (w_0293_, w_1042_, w_1493_);
and (w_1608_, new_in5[6], w_1794_);
nand (w_0275_, w_1250_, w_1329_);
nand (w_2272_, w_1563_, w_1331_);
nand (w_1704_, w_1021_, w_0795_);
nand (w_0568_, new_in23[3], new_in6[3]);
xor (w_2170_, w_0398_, w_0119_);
xor (w_0628_, w_0310_, w_0683_);
or (new_out16[2], w_2238_, w_2294_);
nand (w_0232_, new_in18[2], new_in20[3]);
or (w_0865_, new_in19[0], new_in19[1]);
not (w_0529_, w_0652_);
nand (new_out17[1], w_0452_, w_1536_);
or (w_1923_, w_0793_, w_0337_);
xor (w_0906_, new_in16[2], w_0733_);
nand (w_1643_, w_1792_, w_1227_);
or (w_1168_, w_1926_, w_0850_);
nand (w_0880_, w_0819_, w_0174_);
nand (w_0165_, w_1837_, w_0635_);
xor (w_1268_, new_in21[4], new_in3[4]);
nand (w_0882_, new_in21[2], new_in3[2]);
nand (w_1484_, w_0923_, w_0394_);
xor (w_1732_, new_in20[6], w_0599_);
nand (w_1283_, w_2322_, w_2159_);
xor (w_2225_, w_2047_, w_1222_);
nand (w_1103_, w_1039_, w_1833_);
xor (w_0051_, new_in22[4], w_1440_);
nand (w_0497_, new_in13[3], new_in24[3]);
xor (w_0097_, w_0676_, w_0272_);
nand (w_2239_, w_0695_, new_in12[3]);
nand (w_1341_, new_in5[6], w_0274_);
and (w_1949_, w_0263_, w_2033_);
xor (w_2161_, new_in23[4], w_0854_);
not (w_0313_, w_0800_);
nand (w_2166_, w_2114_, w_2126_);
nand (w_0966_, w_0288_, w_2276_);
and (new_out10[0], w_0375_, w_1862_);
nand (w_0913_, w_0830_, w_0377_);
nand (w_0215_, new_in20[0], w_0348_);
xor (w_1040_, w_1728_, w_2147_);
nand (w_0056_, w_1312_, w_2321_);
xor (w_2042_, new_in5[1], w_1487_);
xor (w_0282_, w_2293_, w_1790_);
nand (w_2031_, w_1905_, w_1737_);
nand (w_0894_, w_0518_, w_0221_);
nand (w_1070_, w_0989_, w_1279_);
nand (w_1447_, new_in9[0], w_0247_);
xor (w_0477_, w_1776_, w_0941_);
xor (w_2126_, w_2274_, w_2188_);
nand (w_1192_, w_1108_, w_0123_);
or (w_2017_, w_0126_, w_0809_);
xor (w_1010_, new_in22[2], new_in21[2]);
and (w_0509_, w_1231_, w_0380_);
xor (w_1497_, w_0075_, w_2185_);
nand (w_1191_, w_0996_, w_1480_);
nand (w_0630_, w_0752_, new_in17[4]);
nand (w_1196_, new_in17[3], new_in10[3]);
xor (w_0054_, new_in18[3], new_in20[4]);
xor (w_1140_, w_1114_, w_2228_);
xor (w_0153_, w_0559_, w_1019_);
or (w_0032_, w_0616_, w_0422_);
nand (w_0356_, w_1905_, w_1541_);
and (w_1602_, w_1625_, w_0745_);
xor (w_2311_, w_0501_, w_2128_);
nand (w_1431_, w_0148_, w_0872_);
and (w_2114_, w_1265_, w_2118_);
xor (w_1869_, w_1826_, w_1633_);
nand (w_0075_, w_0147_, w_0494_);
xor (w_0481_, new_in3[5], w_1729_);
nand (w_0446_, w_1380_, w_0435_);
or (w_0117_, w_1231_, w_1777_);
xor (w_1599_, new_in1[3], new_in9[3]);
nand (w_1760_, w_2300_, w_1174_);
nand (w_1712_, w_0592_, w_0686_);
nand (w_1648_, w_1824_, w_0448_);
nand (w_1101_, w_0263_, w_0018_);
xor (w_1155_, w_2135_, w_2039_);
nand (w_1926_, w_1165_, w_0148_);
and (w_0758_, w_1336_, w_1002_);
xor (w_1569_, w_1315_, w_1107_);
xor (w_2155_, new_in24[2], new_in2[2]);
and (w_0187_, w_1231_, w_1129_);
or (w_2187_, w_0422_, w_1476_);
xor (w_1933_, new_in12[0], new_in12[1]);
or (w_1221_, w_1370_, w_1359_);
nand (w_0721_, w_0025_, w_0093_);
xor (w_1141_, w_1405_, w_0564_);
xor (w_1592_, new_in4[1], w_0860_);
xor (w_2104_, new_in9[0], new_in22[3]);
or (w_1969_, w_0707_, w_0734_);
xor (w_1132_, w_0224_, w_1040_);
and (w_1612_, w_2093_, w_1669_);
and (w_0878_, w_0263_, w_0363_);
nand (w_0513_, new_in10[8], w_1661_);
xor (w_2097_, new_in13[1], new_in13[2]);
xor (w_2056_, w_0324_, w_0479_);
xor (w_0478_, w_2153_, w_1352_);
and (w_1253_, w_1750_, w_1337_);
nand (new_out10[5], w_1449_, w_1406_);
nor (new_out18[3], w_0505_, w_0919_);
nand (w_1675_, w_2038_, w_0349_);
nand (w_0646_, new_in10[8], w_1553_);
and (w_1182_, new_in16[7], w_0011_);
nand (w_1895_, w_0407_, w_2069_);
xor (w_1498_, w_0871_, w_1011_);
nand (w_1402_, new_in10[8], w_1664_);
nand (w_0303_, w_1867_, w_1037_);
nand (w_0672_, new_in10[8], w_1523_);
or (w_1964_, w_1051_, w_1069_);
xor (w_2318_, w_1739_, w_1644_);
xor (w_0708_, w_0526_, w_2320_);
not (w_1161_, new_in12[0]);
xor (w_1208_, new_in8[1], w_0994_);
nand (w_0641_, w_2029_, w_0946_);
nand (w_1480_, w_1289_, w_1367_);
nand (w_1702_, new_in24[4], new_in2[4]);
nand (w_1886_, new_in24[1], new_in2[1]);
nand (w_0535_, w_0619_, w_1861_);
nand (w_2077_, w_2068_, new_in12[2]);
nand (w_0808_, new_in17[2], new_in10[3]);
xor (w_0571_, new_in22[2], new_in14[1]);
nand (w_0786_, new_in16[7], w_0066_);
nand (w_2045_, w_0334_, w_0503_);
and (w_0944_, w_2140_, w_0849_);
nand (w_0709_, w_0084_, w_1351_);
xor (w_1063_, new_in8[4], w_1145_);
not (w_1962_, w_2241_);
or (w_0506_, w_0788_, w_0606_);
and (w_2227_, new_in21[0], new_in3[0]);
nand (w_1148_, w_0869_, w_2230_);
nand (w_0398_, w_0949_, w_1436_);
and (w_1607_, w_0450_, w_0565_);
nor (w_2148_, w_0263_, w_1942_);
and (w_1038_, w_0485_, w_2262_);
or (w_0034_, w_1231_, w_1721_);
or (w_0840_, w_1231_, w_2152_);
xor (w_0955_, w_2273_, w_0214_);
nand (w_1198_, new_in22[2], w_1397_);
nand (w_0121_, w_0017_, w_0387_);
nand (w_0678_, w_1032_, w_0742_);
or (w_2108_, w_1478_, w_1743_);
nand (w_2165_, new_in8[3], w_1461_);
xor (w_1408_, w_1489_, w_2129_);
nand (w_0614_, w_1708_, w_0629_);
or (w_1505_, w_0263_, w_2311_);
xor (w_0066_, w_1666_, w_1542_);
nand (w_0853_, w_0936_, w_1974_);
nand (w_1701_, w_1617_, w_1918_);
nand (w_1396_, w_0428_, w_1443_);
xor (w_1410_, new_in4[3], w_1868_);
xor (w_1565_, new_in5[3], w_0891_);
nand (w_2222_, new_in18[3], new_in20[4]);
xor (w_2142_, w_0188_, w_1951_);
xor (w_0975_, w_2038_, w_0349_);
xor (w_0647_, new_in22[5], new_in9[2]);
or (w_1944_, w_1630_, w_0679_);
xor (w_0002_, w_2229_, w_0360_);
and (w_0399_, w_0597_, w_0502_);
nand (w_0943_, w_1052_, w_2226_);
xor (w_2249_, w_0600_, w_2172_);
or (w_0697_, w_1232_, w_1390_);
nand (w_0182_, new_in22[3], w_1650_);
nand (w_2061_, new_in17[3], new_in10[4]);
nand (w_1212_, w_0613_, w_2265_);
or (w_0692_, w_1193_, w_1592_);
xor (w_2032_, w_0801_, w_0015_);
not (w_1314_, w_1737_);
and (w_1750_, w_0608_, w_0301_);
nand (w_0206_, new_in13[2], new_in24[2]);
xor (w_1735_, new_in7[4], w_0412_);
nand (w_1386_, w_0158_, w_1417_);
nand (w_0098_, new_in20[5], w_1623_);
and (w_1355_, w_0620_, w_0275_);
xor (w_0851_, w_0832_, w_1569_);
nand (w_1200_, w_1677_, w_0470_);
nand (w_1935_, w_0094_, w_1606_);
and (w_1186_, new_in5[6], w_0425_);
xor (w_1778_, w_0162_, w_0466_);
nand (w_1636_, w_1327_, w_0763_);
nand (w_0573_, w_1171_, w_0197_);
and (w_1275_, w_0714_, w_1070_);
and (w_0396_, w_1237_, w_0386_);
nand (w_1459_, w_2251_, w_0424_);
nand (w_1243_, new_in19[2], new_in12[2]);
nand (w_1057_, w_0539_, w_0935_);
nand (w_0597_, new_in5[6], w_1496_);
nand (w_0991_, new_in7[4], new_in8[5]);
nand (new_out8[1], w_1228_, w_1659_);
xor (w_2215_, w_1874_, w_2253_);
xor (w_1310_, w_1956_, w_2192_);
xor (w_2073_, w_1362_, w_0490_);
nand (w_0456_, w_1958_, w_2125_);
nand (w_1867_, w_0923_, w_1321_);
and (new_out9[3], w_0866_, w_0302_);
xor (w_0095_, new_in22[4], new_in21[4]);
and (w_2196_, new_in8[0], new_in1[1]);
and (w_0063_, new_in6[0], new_in11[0]);
nand (w_0766_, w_1568_, w_0550_);
nand (w_1966_, new_in5[5], w_0708_);
xor (w_0501_, w_0458_, w_1343_);
nand (w_1230_, new_in18[2], new_in6[3]);
xor (w_1922_, new_in6[0], new_in18[0]);
nand (w_0163_, w_1486_, w_1879_);
xor (w_1548_, w_1307_, w_0807_);
nand (w_1900_, w_2113_, w_1979_);
nor (w_0170_, w_0263_, w_1555_);
xor (w_0376_, new_in7[1], new_in14[1]);
or (w_1115_, w_1231_, w_1933_);
nand (w_0836_, w_2058_, w_0316_);
nand (w_1536_, w_1892_, w_1213_);
or (w_0566_, w_2093_, w_0361_);
and (w_2071_, w_1519_, w_2157_);
xor (w_0665_, new_in9[5], new_in15[5]);
xor (w_1265_, new_in8[0], new_in1[1]);
nand (w_2184_, new_in12[0], new_in19[0]);
and (new_out15[0], w_1124_, w_1540_);
nor (w_1358_, w_0263_, w_2248_);
or (w_0582_, w_0422_, w_0838_);
nand (w_2265_, w_1863_, w_0823_);
nor (new_out14[4], w_1259_, w_0326_);
nand (w_1956_, w_0189_, w_0312_);
nand (w_0438_, new_in16[7], w_0220_);
nand (w_0299_, w_0351_, w_1910_);
xor (w_2022_, new_in14[0], new_in21[0]);
xor (w_1598_, w_1680_, w_0663_);
nand (w_1628_, w_2280_, w_0257_);
nand (w_0545_, w_0797_, w_1176_);
and (w_0960_, w_1917_, w_1720_);
not (w_1270_, w_1327_);
nand (w_1258_, new_in22[3], new_in16[3]);
nand (w_1491_, w_2206_, w_2170_);
and (w_1757_, w_1231_, w_1714_);
and (new_out16[0], w_2093_, w_1087_);
nand (w_1250_, w_0578_, w_1199_);
nand (w_0374_, w_0967_, w_0496_);
or (w_0252_, w_0338_, w_0480_);
nand (w_2220_, new_in1[2], new_in9[2]);
and (w_2289_, w_1231_, w_0019_);
nand (w_0410_, w_0772_, w_0343_);
nand (w_1908_, w_1231_, w_0078_);
xor (w_1084_, w_0541_, w_1719_);
nand (w_1870_, w_1012_, w_0604_);
xor (w_1350_, w_0673_, w_1871_);
nand (w_1345_, w_1105_, w_0253_);
nand (w_2070_, w_2222_, w_0896_);
nand (w_0869_, w_1396_, w_0153_);
nand (w_1981_, new_in5[6], w_2305_);
nand (w_1997_, w_0376_, w_0881_);
nand (w_0464_, new_in21[4], new_in20[5]);
nand (w_2251_, new_in16[7], w_0622_);
xor (w_0214_, new_in22[2], w_1202_);
nor (w_1433_, w_1647_, new_in17[5]);
xor (w_0171_, w_1457_, w_0000_);
nand (w_1025_, w_0557_, w_0804_);
nand (w_1185_, w_1905_, w_0916_);
nand (w_0129_, w_0907_, w_0156_);
xor (w_1022_, new_in21[2], new_in20[3]);
xor (w_1308_, new_in23[6], w_1693_);
xor (w_1768_, w_0188_, w_1604_);
nand (w_1510_, new_in16[7], w_1823_);
nand (new_out12[0], w_0117_, w_1432_);
xor (w_1097_, new_in21[4], w_2303_);
nand (w_0141_, new_in24[3], new_in2[3]);
nand (new_out11[0], w_2251_, w_1324_);
xor (w_2295_, new_in20[0], w_0861_);
xor (w_0763_, new_in19[4], new_in12[4]);
nand (w_1562_, w_0291_, w_0455_);
nand (w_1642_, new_in22[0], w_1343_);
xor (w_0918_, w_0953_, w_0677_);
and (w_0868_, w_1231_, w_1529_);
xor (w_1769_, new_in12[0], new_in22[0]);
nand (w_0920_, w_2249_, w_1078_);
nand (w_0261_, new_in16[7], w_1797_);
xor (w_1544_, w_1289_, w_1367_);
nand (w_0257_, w_1412_, w_1034_);
xor (w_0916_, w_0966_, w_1720_);
nand (w_2317_, w_0526_, w_2320_);
nand (w_1718_, new_in12[4], new_in15[2]);
xor (w_1249_, new_in14[4], new_in21[4]);
nand (w_0124_, w_2199_, w_1691_);
xor (w_0543_, new_in9[6], new_in1[6]);
nand (w_1420_, new_in4[3], new_in3[3]);
and (new_out3[1], w_0415_, w_0389_);
nand (w_0911_, w_2182_, w_0974_);
nand (w_0307_, new_in21[1], new_in20[2]);
nand (w_1340_, w_1512_, w_1965_);
nand (w_1725_, w_1477_, w_0392_);
xor (w_1458_, w_1312_, w_0313_);
and (w_0357_, new_in19[1], new_in6[0]);
xor (w_0337_, w_1642_, w_2060_);
xor (w_0622_, new_in24[0], new_in2[0]);
nand (w_0634_, new_in5[1], new_in9[2]);
and (new_out1[1], w_1919_, w_1112_);
xor (w_0226_, w_2179_, w_0848_);
nand (w_1122_, w_1587_, w_0185_);
xor (w_1816_, new_in19[5], new_in6[4]);
and (w_1852_, w_1905_, w_1490_);
nand (w_1762_, w_1403_, w_1451_);
xor (w_0698_, new_in5[2], w_1469_);
nand (w_0522_, w_2264_, w_1621_);
nand (w_2098_, w_1072_, w_1608_);
and (w_0608_, new_in7[0], new_in7[1]);
xor (w_1113_, new_in7[5], w_0900_);
xor (w_0821_, new_in21[1], new_in20[2]);
or (w_2218_, w_0422_, w_1571_);
not (w_1766_, new_in23[1]);
nand (w_2260_, w_0250_, w_0548_);
and (w_2028_, new_in10[8], w_2053_);
xor (w_0149_, new_in13[6], new_in24[6]);
xor (w_2085_, w_1116_, w_2186_);
nand (w_1804_, new_in5[6], w_1736_);
and (w_2130_, new_in19[0], w_0022_);
and (w_0804_, new_in16[7], w_1985_);
nand (new_out12[6], w_1856_, w_0243_);
and (w_1284_, w_2239_, w_0815_);
xor (w_1546_, w_0912_, w_1338_);
xor (w_1633_, new_in23[5], new_in6[5]);
or (w_0979_, w_2093_, w_0775_);
nand (w_1055_, w_0560_, w_0791_);
or (w_2304_, w_2093_, w_0737_);
xor (w_2321_, w_1209_, w_2120_);
and (w_2206_, w_2084_, w_1812_);
or (w_0627_, new_in13[2], new_in13[4]);
nand (w_1335_, new_in5[6], new_in5[0]);
xor (w_1187_, new_in1[2], new_in9[2]);
nand (w_2047_, w_0547_, w_1055_);
xor (w_1088_, w_0485_, w_2262_);
or (w_0504_, new_in8[2], w_0086_);
xor (w_1720_, w_0852_, w_0289_);
and (w_1166_, new_in5[6], w_1276_);
nand (w_0956_, w_0642_, w_1509_);
nand (w_0969_, new_in5[4], w_0628_);
xor (w_2281_, new_in23[1], new_in6[1]);
or (w_1240_, w_1575_, w_1541_);
nand (w_2291_, new_in18[5], new_in11[5]);
and (w_0240_, new_in3[0], w_0128_);
nand (w_1531_, w_0075_, w_1524_);
xor (w_0069_, w_0383_, w_1938_);
xor (w_0359_, new_in18[1], new_in11[1]);
nand (w_1273_, w_1234_, w_1745_);
nand (w_1837_, new_in11[1], w_0143_);
nand (w_1551_, new_in10[8], w_0489_);
xor (w_0687_, w_1380_, w_0435_);
nand (w_0318_, w_1713_, w_2025_);
xor (w_0242_, w_1270_, w_0763_);
xor (w_0904_, new_in4[3], new_in3[3]);
not (w_2137_, new_in22[5]);
nand (w_0922_, w_1320_, w_1772_);
or (w_2275_, w_2273_, w_0214_);
xor (w_1469_, w_2097_, w_1511_);
nand (w_0332_, new_in18[1], new_in6[2]);
nand (w_2277_, w_0871_, w_1011_);
and (w_0403_, w_1231_, w_0065_);
nand (w_1756_, w_0263_, w_0124_);
nand (w_0074_, w_1819_, w_0178_);
nand (new_out9[5], w_0048_, w_1130_);
nand (w_1425_, new_in4[2], w_0445_);
nand (w_0613_, w_1011_, w_0549_);
nand (w_1994_, w_1849_, w_0818_);
xor (w_0828_, new_in13[3], new_in24[3]);
xor (w_0479_, w_0164_, w_2181_);
and (w_0010_, new_in16[7], w_0577_);
nand (w_1073_, w_1234_, w_0229_);
and (w_2129_, w_1993_, w_0777_);
or (w_0236_, w_1820_, w_0009_);
and (w_2099_, w_1777_, w_1818_);
nand (w_1825_, new_in5[6], w_0352_);
xor (w_2147_, w_1486_, w_1879_);
nand (w_1875_, w_1629_, w_2014_);
xor (w_1541_, w_1372_, w_0443_);
nand (w_1843_, new_in3[4], w_1544_);
xor (w_1806_, w_0457_, w_0689_);
nand (w_0184_, w_1231_, w_0159_);
xor (w_0060_, new_in22[4], new_in16[4]);
nand (w_0636_, w_1666_, w_0940_);
xor (w_1367_, new_in4[4], new_in2[4]);
nand (w_1815_, w_0947_, w_1064_);
nand (w_1841_, w_1902_, w_1136_);
or (w_1842_, w_0338_, w_1471_);
and (w_0448_, w_0263_, w_0356_);
nand (w_0298_, w_1057_, w_2100_);
nand (w_1545_, new_in18[4], new_in6[5]);
xor (w_2242_, w_1747_, w_1120_);
nand (w_0802_, w_0567_, w_2281_);
xor (w_0783_, new_in4[2], w_0445_);
xor (w_1942_, w_2219_, w_1988_);
xor (w_0411_, w_2143_, w_1844_);
or (w_2106_, w_0263_, w_0147_);
nor (w_0412_, w_1446_, new_in7[2]);
and (new_out9[4], w_0770_, w_0271_);
and (w_1931_, new_in10[8], w_0639_);
xor (w_1422_, w_0327_, w_0901_);
nand (w_0617_, w_0697_, w_1570_);
xor (w_1343_, new_in23[0], w_1913_);
xor (w_0901_, w_1728_, w_0700_);
xor (w_1883_, new_in11[1], w_0143_);
nand (new_out13[5], w_1400_, w_1775_);
nor (new_out6[3], w_1346_, w_1513_);
and (w_0623_, w_0136_, w_0886_);
or (w_1755_, w_1232_, w_2308_);
or (w_1174_, w_2255_, w_2034_);
or (w_1519_, w_0772_, w_0343_);
xor (w_0625_, new_in13[5], new_in24[5]);
or (w_2288_, w_0501_, w_2128_);
nand (w_2117_, new_in23[1], new_in6[1]);
nand (w_2183_, w_1601_, w_1510_);
nand (w_0551_, w_2047_, w_1222_);
xor (w_1780_, w_1051_, w_1069_);
xor (w_0838_, w_0632_, w_1210_);
xor (w_0434_, new_in18[0], new_in11[0]);
xor (w_0704_, new_in14[3], new_in22[3]);
nand (w_1377_, w_0336_, w_1661_);
xor (w_1125_, w_0929_, w_2237_);
xor (w_0861_, new_in7[0], new_in14[0]);
or (w_2261_, w_0832_, w_1569_);
nand (w_0003_, new_in7[5], new_in15[5]);
xor (w_2001_, w_0063_, w_1883_);
xor (w_1597_, w_1312_, w_2321_);
and (new_out17[2], w_0487_, w_0767_);
xor (w_1839_, w_0240_, w_2086_);
nand (w_0039_, w_0717_, w_1800_);
or (w_1793_, w_1231_, w_2088_);
xor (w_1797_, w_0590_, w_1602_);
xor (w_1823_, w_2261_, w_0069_);
xor (w_0559_, w_1665_, w_0810_);
xor (w_0038_, w_0288_, w_2276_);
nand (new_out17[6], w_1811_, w_1924_);
and (w_1360_, new_in10[8], w_0515_);
xor (w_0419_, w_1766_, w_0556_);
xor (w_1879_, new_in3[4], w_1544_);
nand (w_0557_, w_2324_, w_1050_);
nand (w_0037_, w_0922_, w_1464_);
or (w_0130_, new_in20[0], w_0348_);
nand (w_0302_, new_in16[7], w_0873_);
and (w_1315_, w_2287_, w_2286_);
nand (w_0656_, w_2162_, w_1221_);
or (w_1754_, w_2093_, w_1980_);
nand (w_1512_, w_2132_, w_0173_);
nand (new_out2[0], w_0117_, w_1254_);
not (w_0644_, w_2171_);
nand (w_0732_, w_1008_, w_0201_);
or (w_1577_, w_1231_, w_1088_);
nand (w_1426_, w_0524_, w_1111_);
and (new_out9[1], w_1505_, w_0728_);
nand (w_0655_, w_0944_, w_1363_);
or (w_1503_, new_in16[7], w_2254_);
and (w_2282_, new_in20[0], w_0861_);
xor (w_0632_, w_0050_, w_0749_);
nand (w_2278_, w_0870_, w_1672_);
nand (w_1972_, w_0173_, w_0794_);
xor (w_0201_, new_in21[3], new_in20[4]);
nand (w_1507_, w_0459_, w_1110_);
and (w_0572_, w_2071_, w_2240_);
or (w_2300_, w_1231_, w_1175_);
nand (new_out14[0], w_2272_, w_1939_);
xor (w_1509_, w_0423_, w_1249_);
xor (w_0941_, new_in19[3], new_in6[2]);
xor (w_0235_, w_1262_, w_1201_);
or (w_1219_, new_in7[4], w_1252_);
xor (w_1019_, w_0120_, w_1288_);
nand (w_0449_, w_0184_, w_0963_);
nand (w_1033_, w_0572_, w_1850_);
and (w_2144_, new_in13[0], new_in1[0]);
nand (w_0554_, w_1016_, w_0889_);
nand (w_0717_, w_1973_, w_1898_);
nand (w_0092_, new_in20[2], w_0975_);
and (new_out15[1], w_0339_, w_1077_);
nand (w_2241_, w_1888_, w_1704_);
nand (w_1456_, new_in14[4], new_in22[5]);
nand (w_1506_, w_1091_, w_0519_);
nand (w_1379_, w_0263_, w_1762_);
nand (w_1373_, new_in17[4], new_in10[4]);
nand (w_2072_, new_in22[2], w_2104_);
nand (w_0291_, w_0923_, w_1934_);
and (w_1820_, w_2198_, w_0287_);
xor (w_1737_, w_1394_, w_0533_);
xor (w_0128_, new_in4[0], new_in2[0]);
or (w_1872_, w_1927_, w_0824_);
xor (w_1309_, new_in13[4], new_in5[4]);
xor (w_0373_, w_0067_, w_0042_);
nand (w_0896_, w_2243_, w_0054_);
or (w_0690_, new_in17[3], w_0807_);
xor (w_0229_, w_0518_, w_0221_);
nand (w_1393_, w_0529_, w_0196_);
nand (new_out4[2], w_1220_, w_0254_);
xor (w_0314_, w_1262_, w_0787_);
nand (w_0159_, w_0914_, w_1137_);
nand (w_1758_, new_in21[3], w_2056_);
nand (w_0676_, w_0212_, w_1589_);
nand (w_1158_, new_in3[3], w_1970_);
not (w_0507_, new_in19[1]);
and (w_1414_, w_1226_, w_0392_);
nand (w_1451_, new_in5[6], w_0251_);
nand (w_0363_, w_1905_, w_2306_);
xor (w_2259_, w_0520_, w_0516_);
nand (w_0779_, w_2057_, w_0648_);
nand (w_0335_, w_2219_, w_1988_);
nand (w_0780_, w_2093_, w_0899_);
nand (w_1605_, w_2296_, w_1192_);
xor (w_0793_, new_in22[0], w_1343_);
nand (w_1054_, w_2059_, w_0980_);
nand (w_1356_, w_2314_, w_1963_);
xor (w_0491_, w_1312_, w_0293_);
xor (w_0316_, w_0006_, w_1329_);
nand (w_1387_, new_in11[2], w_0785_);
xor (w_0352_, new_in5[4], w_0806_);
or (w_2141_, new_in18[0], new_in20[1]);
and (w_1689_, new_in24[0], new_in2[0]);
nor (w_1912_, w_1231_, w_1899_);
nand (w_0755_, w_1488_, w_2008_);
nand (w_1532_, w_0960_, w_0242_);
nand (w_2312_, w_1701_, w_0698_);
and (w_2105_, w_2065_, w_1645_);
nand (w_0724_, new_in12[1], w_0376_);
or (w_2036_, w_1642_, w_2060_);
xor (w_1383_, new_in20[5], w_1623_);
xor (w_1901_, new_in19[1], new_in17[1]);
and (w_0079_, w_1488_, w_0161_);
nand (w_0892_, w_0856_, w_1299_);
nor (new_out8[5], w_0659_, w_1893_);
nand (w_1889_, w_0292_, w_1146_);
nand (w_2197_, new_in13[0], w_0250_);
nand (w_1478_, w_1485_, w_0179_);
nand (w_0455_, new_in10[8], w_1013_);
xor (w_0983_, new_in14[6], new_in7[6]);
nand (new_out3[2], w_0780_, w_0961_);
or (w_0029_, w_2093_, w_0097_);
or (w_1936_, w_0800_, w_2057_);
xor (w_2111_, new_in20[4], w_1810_);
nor (w_0202_, w_2295_, w_0268_);
nand (w_1586_, w_1109_, w_2142_);
nand (w_1543_, new_in21[2], new_in20[3]);
or (w_1558_, w_0202_, w_0587_);
nand (w_1864_, w_1194_, w_1782_);
xor (w_1312_, new_in22[2], w_2104_);
nor (w_0659_, w_0263_, w_1225_);
xor (w_0999_, new_in7[1], new_in15[1]);
xor (w_0863_, w_1923_, w_1546_);
xor (w_1965_, w_0293_, w_0699_);
xor (w_1153_, new_in8[3], w_1461_);
xor (w_2122_, new_in19[1], new_in6[0]);
nand (w_1625_, w_0401_, w_0848_);
nand (w_2243_, w_0232_, w_2191_);
nand (w_0530_, w_0585_, w_1947_);
xor (w_1029_, w_0843_, w_1167_);
nand (w_2219_, w_0328_, w_0956_);
not (w_0576_, w_0748_);
and (w_1738_, new_in1[0], new_in9[0]);
not (w_0164_, new_in11[3]);
or (w_0203_, w_1231_, w_1132_);
and (w_0431_, w_0775_, w_1457_);
xor (w_1550_, w_0650_, w_1239_);
xor (w_0220_, new_in12[0], w_0861_);
or (w_1539_, new_in19[2], w_0865_);
nand (w_0694_, w_0241_, w_0641_);
nand (w_0025_, w_1699_, w_1264_);
and (w_1452_, new_in18[0], new_in11[0]);
nand (w_1977_, new_in5[2], w_1469_);
nand (w_0971_, w_1325_, w_2139_);
xor (w_0917_, new_in22[0], w_0244_);
xor (w_1604_, w_2092_, w_0661_);
nand (w_0450_, new_in1[3], new_in8[2]);
xor (w_0683_, w_0837_, w_1911_);
nand (w_1809_, w_1042_, w_1493_);
nand (w_2292_, w_1905_, w_0653_);
nand (w_2092_, w_1715_, w_0322_);
nand (w_0771_, w_1649_, w_1517_);
nand (w_0816_, new_in8[2], w_0086_);
nand (w_0825_, w_1997_, w_1364_);
and (w_0929_, w_1955_, w_0932_);
or (w_1857_, w_1139_, w_0259_);
and (w_0498_, w_1859_, w_0868_);
xor (w_1417_, new_in12[1], new_in22[1]);
nand (w_0462_, w_0293_, w_0699_);
nand (new_out6[1], w_1793_, w_2201_);
xor (w_0133_, new_in5[2], new_in13[2]);
nand (w_1619_, w_1038_, w_1881_);
and (w_1928_, w_1922_, w_0542_);
nand (w_1392_, w_2043_, w_1138_);
xor (w_1728_, w_1753_, w_0137_);
nand (w_1313_, w_0456_, w_1774_);
xor (w_0435_, new_in7[4], new_in8[5]);
nand (w_1660_, w_0400_, w_1786_);
and (w_0519_, w_1234_, w_0045_);
xor (w_1218_, w_1849_, w_1027_);
nand (w_2209_, w_0681_, w_1654_);
nand (w_1131_, w_0126_, w_1184_);
nand (w_0635_, w_0063_, w_1883_);
nand (w_1444_, new_in4[3], w_1868_);
nand (w_1302_, new_in5[6], w_0105_);
nand (w_1649_, new_in1[2], new_in13[2]);
nand (w_1000_, w_2168_, new_in17[3]);
nand (w_1449_, w_1231_, w_1450_);
nand (w_0353_, w_1905_, w_1945_);
nand (w_1096_, w_0973_, w_1418_);
nand (w_0276_, w_2235_, w_1022_);
xor (w_1173_, new_in13[5], new_in1[5]);
nand (w_0026_, w_0874_, w_1609_);
nand (w_2037_, w_0871_, w_0392_);
and (w_0250_, w_2093_, new_in5[6]);
or (w_0469_, w_1283_, w_1768_);
nand (w_1332_, new_in20[1], w_0982_);
and (w_0517_, w_1114_, w_2228_);
xor (w_2248_, w_1376_, w_1348_);
xor (w_2163_, w_2105_, w_0401_);
and (w_0457_, new_in22[0], w_0244_);
nand (w_0619_, new_in16[4], w_2161_);
nand (new_out16[1], w_0285_, w_0102_);
nand (w_2263_, w_2285_, w_0744_);
not (w_0260_, w_0094_);
nand (w_0428_, w_2048_, w_2208_);
or (w_1026_, w_1232_, w_1769_);
nand (w_1783_, w_1975_, w_1291_);
nand (w_2096_, new_in5[6], w_1438_);
or (w_0932_, w_1717_, w_0140_);
xor (w_0592_, new_in17[4], new_in10[4]);
nand (w_0768_, new_in1[5], new_in9[5]);
not (w_1634_, new_in13[4]);
nand (w_1204_, new_in7[2], new_in8[3]);
xor (w_0935_, w_0881_, w_1004_);
nand (w_0297_, new_in4[1], new_in3[1]);
and (new_out12[4], w_1577_, w_0440_);
xor (w_2048_, w_1152_, w_0736_);
xor (w_1288_, new_in13[4], new_in24[4]);
xor (w_2169_, w_1694_, w_0722_);
nand (w_0620_, new_in16[4], w_2147_);
nand (w_0642_, w_0779_, w_0465_);
nand (w_0134_, w_1766_, new_in12[1]);
nand (w_2064_, new_in3[5], w_1729_);
or (w_0045_, w_0228_, w_0150_);
nand (w_0742_, w_1927_, w_0824_);
xor (w_1256_, w_0122_, w_1796_);
nand (w_2274_, w_1882_, w_2302_);
nand (w_1299_, w_0340_, w_0194_);
nand (w_0484_, w_1191_, w_0976_);
nand (w_2025_, w_1394_, w_0533_);
and (new_out7[0], w_1707_, w_0371_);
nand (w_1432_, w_1231_, w_2005_);
xor (w_2054_, w_1095_, w_1153_);
and (w_1744_, new_in4[0], new_in2[0]);
nand (w_1937_, w_1905_, w_0962_);
nand (new_out11[6], w_1409_, w_1179_);
nor (w_1887_, w_1231_, w_0397_);
nand (w_0440_, w_0341_, w_1757_);
and (w_1242_, w_1420_, w_0073_);
nand (w_0091_, w_0263_, new_in5[6]);
nand (w_0930_, w_1361_, w_0135_);
and (w_0267_, new_in8[0], w_1467_);
xor (w_0101_, new_in11[5], w_0525_);
xor (w_0119_, w_0700_, w_0423_);
nand (w_0452_, w_0731_, w_0421_);
xor (w_1238_, w_1426_, w_1295_);
and (w_2186_, w_1813_, w_0134_);
nand (w_0544_, new_in16[7], w_0803_);
nand (w_1042_, w_1255_, w_0037_);
nand (w_2195_, w_1319_, w_2062_);
nand (w_1578_, w_0052_, w_0490_);
xor (w_2118_, w_2196_, w_1119_);
xor (w_1348_, new_in22[3], new_in21[3]);
and (w_1411_, new_in5[6], w_1168_);
nand (w_0345_, new_in13[1], new_in1[1]);
nand (w_0106_, w_2093_, w_0530_);
nand (w_2107_, w_0610_, w_0108_);
nand (w_0673_, w_1456_, w_0573_);
nand (w_2087_, w_1231_, w_1580_);
nand (w_2235_, w_0307_, w_1160_);
or (w_0842_, w_1211_, w_0040_);
nand (w_0939_, w_2295_, w_0268_);
and (w_2124_, w_2127_, w_1354_);
nand (w_1915_, new_in4[2], new_in3[2]);
nand (w_0127_, new_in5[6], w_1067_);
nand (w_1139_, w_0468_, w_0058_);
xor (w_0194_, new_in21[2], w_0343_);
xor (w_2315_, new_in7[1], new_in8[2]);
xor (w_1751_, new_in5[3], new_in13[3]);
or (w_2214_, w_1231_, w_1516_);
xor (w_1868_, w_1205_, w_0512_);
xor (w_0067_, w_0499_, w_0665_);
nand (w_1276_, w_0517_, w_0133_);
nand (w_1772_, w_0240_, w_2086_);
xor (w_1516_, w_1109_, w_2142_);
nand (w_2133_, new_in5[6], w_0024_);
xor (w_2101_, w_0429_, w_2063_);
nand (w_0044_, new_in16[7], w_2216_);
nand (w_1761_, w_1189_, w_1597_);
or (w_0803_, w_1522_, w_1310_);
or (w_0160_, w_2093_, w_0583_);
xor (w_0112_, w_2317_, w_0918_);
and (w_0764_, w_0827_, w_1375_);
nand (w_0245_, new_in16[7], w_1195_);
and (w_1007_, w_1231_, w_1026_);
nand (new_out13[1], w_0595_, w_0618_);
nand (w_0788_, w_1389_, w_0334_);
xor (w_2060_, new_in22[1], w_0419_);
nand (w_0019_, w_0522_, w_0085_);
nand (w_0928_, w_2018_, w_0187_);
xor (w_1954_, w_0729_, w_1280_);
and (new_out11[5], w_0985_, w_0598_);
xor (w_0677_, new_in13[6], w_1408_);
nand (w_0028_, w_0263_, w_0449_);
or (w_2008_, new_in16[3], w_1650_);
or (w_1745_, w_2127_, w_1354_);
xor (w_0546_, new_in22[1], new_in21[1]);
xor (w_0611_, w_0205_, w_0478_);
or (w_0948_, w_1231_, w_1550_);
nand (w_1835_, new_in4[2], new_in2[2]);
nand (w_1205_, w_0141_, w_1535_);
nand (w_2006_, new_in21[3], new_in3[3]);
or (w_1903_, w_1575_, w_0903_);
and (w_1655_, w_0263_, w_1799_);
and (w_0743_, w_1161_, new_in23[0]);
xor (w_1818_, w_1180_, w_0999_);
xor (w_0660_, w_1925_, w_0070_);
nor (new_out5[4], w_1445_, w_0498_);
and (w_0777_, new_in13[3], w_0627_);
xor (w_1974_, new_in5[4], w_0628_);
nand (w_0224_, w_1640_, w_0071_);
nand (w_1254_, w_0926_, w_0473_);
nand (w_0870_, w_1230_, w_1895_);
and (w_2293_, w_0431_, w_1588_);
nand (w_0062_, w_0074_, w_1684_);
and (w_1277_, w_2093_, w_1773_);
xor (w_1877_, w_0950_, w_1005_);
xor (w_2039_, w_0401_, w_1951_);
xor (w_0981_, w_2263_, w_0855_);
nand (w_0651_, w_0263_, w_1573_);
and (w_1764_, w_1231_, w_2158_);
xor (w_0658_, new_in4[0], w_2190_);
nand (w_0831_, new_in5[6], w_2076_);
xor (w_0185_, new_in12[5], new_in15[3]);
xor (w_2276_, w_0576_, w_1521_);
or (w_1448_, w_0422_, w_0790_);
nand (w_1248_, w_1724_, w_0372_);
and (w_0473_, w_1231_, w_1098_);
and (w_0476_, w_1231_, w_1506_);
nand (w_1035_, w_1236_, w_2278_);
nand (w_2102_, w_1917_, w_1720_);
nand (w_1596_, w_2006_, w_0193_);
xor (w_2038_, new_in17[2], new_in10[2]);
and (w_0889_, new_in5[6], w_1878_);
nand (w_1465_, w_1312_, w_0800_);
nand (w_1143_, w_1231_, w_1374_);
or (w_0718_, w_2243_, w_0054_);
not (w_0695_, new_in23[3]);
xor (w_1316_, new_in5[3], w_1695_);
nand (w_2217_, w_1457_, w_0000_);
not (w_0710_, new_in22[3]);
nand (w_1428_, w_0747_, w_0869_);
xor (w_0305_, w_0572_, w_1850_);
or (w_2174_, w_0713_, w_0670_);
and (w_0607_, new_in16[7], w_1395_);
nand (w_0681_, w_1283_, w_1768_);
xor (w_0256_, w_1967_, w_0223_);
and (w_0087_, w_1231_, w_0674_);
xor (w_2171_, new_in19[5], new_in17[5]);
nand (w_1587_, w_1718_, w_0062_);
xor (w_0867_, w_0649_, w_1309_);
nand (new_out7[4], w_0280_, w_1594_);
and (w_1814_, new_in13[0], new_in5[0]);
xor (w_0626_, new_in24[3], new_in2[3]);
nand (w_2302_, w_2196_, w_1119_);
and (w_2294_, w_2093_, w_1635_);
nand (w_1320_, new_in3[1], w_0811_);
nand (w_0253_, new_in16[7], w_1104_);
or (w_2035_, w_0263_, w_0793_);
nand (w_1117_, w_2074_, w_1302_);
or (w_0818_, new_in17[5], new_in10[5]);
xor (w_1015_, w_2233_, w_0925_);
nand (w_0499_, w_0001_, w_2247_);
xor (w_1752_, new_in23[1], new_in12[1]);
or (w_1662_, w_0508_, w_0294_);
xor (w_1650_, new_in23[3], w_1548_);
nand (w_1860_, w_0775_, w_2016_);
and (w_0207_, w_0945_, w_0681_);
and (w_0218_, new_in1[1], w_1663_);
xor (w_1106_, w_0989_, w_1279_);
nand (w_1409_, w_0263_, w_1117_);
xor (w_1247_, w_0884_, w_0411_);
xor (w_1397_, new_in23[2], w_1560_);
nand (w_1455_, w_0464_, w_2049_);
nand (w_0515_, w_1502_, w_2256_);
nand (new_out4[5], w_0072_, w_1434_);
or (w_0601_, new_in5[0], new_in5[1]);
nand (w_1051_, w_0883_, w_1141_);
nand (w_0368_, w_2277_, w_1246_);
xor (w_0301_, new_in7[2], new_in7[1]);
nand (w_0217_, w_0125_, w_1593_);
xor (w_0976_, new_in4[5], new_in2[5]);
xor (w_0070_, new_in22[1], w_0376_);
nand (w_1631_, w_2179_, w_0042_);
nand (w_0391_, new_in10[8], w_0282_);
nand (w_1001_, new_in19[3], w_0690_);
xor (w_2257_, new_in4[2], new_in2[2]);
nand (new_out14[5], w_0774_, w_0329_);
nand (w_2013_, new_in13[1], new_in13[2]);
or (w_0408_, w_1231_, w_1876_);
or (w_0729_, w_1747_, w_1120_);
xor (w_1014_, w_1607_, w_0540_);
and (w_1003_, w_1231_, w_0979_);
nand (w_0216_, new_in17[3], w_0807_);
nand (w_2074_, w_1905_, w_1015_);
xor (w_2228_, new_in5[1], new_in13[1]);
nand (w_0754_, w_1234_, w_0746_);
xor (w_1089_, w_2108_, w_1269_);
xor (w_1585_, w_0710_, w_1650_);
nand (w_2223_, w_2140_, w_1186_);
nand (w_1043_, w_1452_, w_0359_);
xor (w_1891_, new_in20[1], w_0982_);
xor (w_0689_, new_in22[1], w_1839_);
nand (w_1620_, w_1918_, w_0169_);
nand (w_0080_, w_0978_, w_1437_);
or (w_0198_, w_2314_, w_1402_);
or (w_1986_, new_in12[0], new_in19[0]);
not (w_0852_, w_0333_);
nand (w_2132_, w_1202_, w_2259_);
nand (w_1652_, w_2093_, w_0100_);
nand (w_0927_, w_1231_, w_1562_);
nand (w_1742_, w_2223_, w_1248_);
nand (w_1775_, new_in5[6], w_1626_);
and (w_0377_, w_0923_, w_1240_);
nand (w_0076_, w_0482_, w_1748_);
xor (w_2078_, w_0099_, w_0101_);
xor (w_1790_, new_in18[5], new_in11[5]);
nand (w_0152_, w_1103_, w_1187_);
xor (w_0199_, new_in23[5], w_1638_);
xor (w_1661_, w_0026_, w_1765_);
nor (new_out5[2], w_1887_, w_1916_);
nand (w_2164_, w_0457_, w_0689_);
xor (w_0269_, new_in1[4], new_in8[4]);
nand (new_out2[4], w_1044_, w_0968_);
and (w_2314_, new_in21[0], w_1960_);
nand (w_2310_, w_0353_, w_0315_);
xor (w_1988_, w_2179_, w_1123_);
nand (w_2082_, new_in5[6], w_0041_);
nand (new_out14[3], w_1233_, w_1622_);
nand (w_1733_, new_in9[2], new_in15[2]);
or (w_0910_, w_0091_, w_1265_);
nand (w_0801_, w_2066_, w_0563_);
or (w_0986_, new_in16[3], w_0293_);
xor (w_1802_, new_in20[0], w_2022_);
nand (w_1289_, w_2080_, w_1056_);
not (w_1477_, new_in22[2]);
nand (w_1710_, w_1311_, w_1097_);
nand (w_1215_, w_1092_, w_1727_);
nand (new_out16[3], w_0270_, w_0103_);
nand (w_0770_, w_0495_, w_0239_);
xor (w_1726_, w_1212_, w_1404_);
nand (w_2081_, w_0248_, w_1646_);
nand (w_0354_, w_2210_, w_1840_);
nand (w_1362_, w_0796_, w_1546_);
and (w_0324_, w_1387_, w_0586_);
nand (w_0555_, w_0224_, w_1040_);
and (w_1989_, w_2007_, w_1126_);
and (w_0209_, new_in23[3], new_in12[3]);
xor (w_0480_, w_0126_, w_0809_);
not (w_2168_, new_in19[3]);
nand (w_1991_, w_1564_, w_0971_);
xor (w_1553_, w_0775_, w_1457_);
xor (w_0196_, w_1839_, w_1920_);
or (w_2245_, new_in8[0], w_1705_);
and (w_0953_, w_1047_, w_2301_);
nand (w_1323_, w_1231_, w_0645_);
nand (w_0900_, w_1219_, w_0562_);
xor (w_0871_, new_in7[2], new_in14[2]);
and (w_0081_, w_1306_, w_0266_);
and (w_0843_, w_0402_, w_0233_);
xor (w_1920_, w_2227_, w_2041_);
xor (w_1036_, new_in1[2], new_in8[2]);
not (w_0022_, new_in17[0]);
nand (w_2011_, new_in16[7], w_2190_);
nor (w_1992_, w_1231_, w_0915_);
xor (w_1464_, new_in3[2], w_1549_);
and (w_1291_, w_0263_, w_1147_);
xor (w_1638_, w_0644_, w_1108_);
not (w_1671_, w_1103_);
nand (w_0534_, w_1977_, w_2312_);
nand (w_1162_, w_2067_, w_0828_);
nor (w_1445_, w_1231_, w_2319_);
nand (w_1327_, w_2046_, w_2023_);
xor (w_0413_, w_0267_, w_1208_);
and (w_0680_, w_2323_, w_0016_);
nand (w_0537_, w_1260_, w_1339_);
xor (w_0360_, w_2137_, new_in21[5]);
nand (w_1489_, new_in13[5], w_1634_);
xor (w_1727_, new_in19[1], new_in12[1]);
and (w_1828_, new_in12[0], w_0861_);
xor (w_0150_, new_in17[3], new_in10[3]);
nand (w_0407_, w_0332_, w_2177_);
xor (w_0881_, new_in21[0], new_in20[1]);
nand (w_0379_, w_1071_, w_0269_);
xor (w_1731_, w_0426_, w_2315_);
and (w_0958_, w_0773_, w_1238_);
and (w_1298_, w_1905_, w_0418_);
xor (w_0800_, new_in7[3], new_in14[3]);
nand (w_0968_, new_in5[6], w_2299_);
nand (w_2200_, w_0923_, w_2194_);
and (w_1384_, new_in19[0], new_in17[0]);
xor (w_0046_, w_1412_, w_1034_);
xor (w_1960_, new_in6[0], new_in11[0]);
and (w_0923_, w_2093_, new_in16[7]);
xor (w_0325_, w_1897_, w_2027_);
and (w_0169_, new_in5[6], w_0213_);
not (w_0772_, w_2001_);
and (w_1827_, w_1231_, w_0646_);
and (w_0560_, new_in17[0], new_in10[1]);
and (w_1376_, w_1846_, w_1010_);
xor (w_2309_, w_0406_, w_1700_);
or (w_1794_, w_1428_, w_0373_);
xor (w_0648_, new_in14[3], new_in21[3]);
nand (w_0973_, w_0308_, w_1852_);
xor (w_2120_, new_in12[3], new_in15[1]);
and (w_1615_, w_0816_, w_0504_);
nand (w_0760_, w_0395_, w_0300_);
nand (w_1753_, w_2156_, w_2072_);
nand (w_0585_, w_0136_, w_1778_);
nand (w_0227_, w_1110_, w_1978_);
and (w_0372_, w_1905_, w_0447_);
nand (w_1979_, w_2241_, w_1534_);
nand (w_0856_, new_in21[2], w_0343_);
xor (w_2088_, new_in5[0], new_in5[1]);
and (w_1206_, w_2165_, w_0654_);
xor (w_2303_, w_0614_, w_1854_);
and (w_0104_, new_in5[6], w_1475_);
nand (w_1124_, w_0263_, w_2081_);
and (w_1226_, new_in12[0], new_in12[1]);
xor (w_1286_, w_1922_, w_0542_);
nand (w_1217_, new_in16[7], w_1030_);
nand (w_2029_, w_0427_, w_1399_);
or (w_1847_, w_0263_, w_1031_);
nand (w_2296_, new_in19[5], new_in17[5]);
nand (w_0096_, w_1326_, w_0559_);
nand (w_0103_, new_in10[8], w_1210_);
and (w_1679_, w_0521_, w_0475_);
nand (w_1973_, new_in7[1], new_in15[1]);
xor (w_0733_, w_2068_, w_1560_);
nand (w_0271_, new_in16[7], w_0664_);
xor (w_1011_, w_0358_, w_0821_);
nand (w_0725_, w_2234_, w_1313_);
nand (w_1694_, w_1685_, w_1583_);
xor (w_2284_, new_in4[5], w_0306_);
nand (w_0909_, new_in18[2], new_in11[2]);
or (w_0084_, w_1033_, w_1317_);
xor (w_0137_, new_in22[4], new_in9[1]);
nand (w_1002_, w_0801_, w_0015_);
nand (w_2229_, w_1334_, w_0095_);
and (w_1027_, w_0451_, w_0818_);
nand (w_1151_, new_in20[2], w_2138_);
nor (w_1259_, w_1231_, w_2054_);
and (w_1834_, w_2293_, w_1790_);
nand (w_1272_, new_in18[1], new_in11[1]);
and (w_0964_, w_1905_, w_1857_);
xor (w_1805_, new_in16[5], w_0188_);
nand (w_0329_, new_in5[6], w_0204_);
nand (w_1785_, new_in4[5], new_in2[5]);
nand (w_0437_, new_in5[3], w_0891_);
xor (w_2019_, w_0668_, w_1657_);
xor (w_1300_, new_in19[6], new_in6[5]);
nand (w_0769_, w_1423_, w_0575_);
xor (w_2152_, new_in5[2], w_0601_);
xor (w_1552_, w_0557_, w_1463_);
not (w_0263_, new_in16[7]);
nand (w_2083_, w_0198_, w_1007_);
and (w_1326_, w_0958_, w_2048_);
nand (new_out18[1], w_0298_, w_0651_);
nand (w_0817_, w_1477_, w_1202_);
nand (w_0071_, w_0030_, w_0491_);
nand (w_1716_, w_0092_, w_1815_);
nand (w_1529_, new_in10[8], w_1789_);
nand (w_1622_, new_in5[6], w_0621_);
nand (w_0116_, w_0263_, w_0219_);
xor (w_1801_, new_in14[3], new_in22[4]);
xor (w_0533_, new_in23[2], new_in6[2]);
nand (w_1924_, new_in10[8], w_1157_);
and (w_1193_, new_in4[0], w_2190_);
or (w_0004_, w_1401_, w_2009_);
xor (w_1467_, new_in7[0], new_in7[1]);
and (w_1821_, w_0263_, w_1046_);
nand (new_out8[6], w_1756_, w_0261_);
nand (w_0595_, w_1231_, w_0080_);
or (w_0180_, w_1231_, w_2318_);
not (w_2154_, w_0771_);
or (w_0115_, w_0517_, w_0133_);
and (w_2269_, new_in5[6], w_1581_);
nand (w_0719_, new_in22[1], w_1839_);
nand (w_1629_, new_in20[4], w_1810_);
nand (w_0461_, w_1231_, w_2183_);
nand (w_1819_, new_in12[3], new_in15[1]);
xor (w_1416_, w_0998_, w_1410_);
nand (w_0048_, w_0263_, w_2211_);
not (w_0367_, new_in13[3]);
nand (w_0812_, w_0896_, w_0706_);
nand (w_0195_, new_in5[6], w_2115_);
or (w_2127_, w_1913_, w_0139_);
xor (w_1993_, new_in13[5], new_in13[4]);
xor (w_1415_, new_in11[6], w_2244_);
nand (w_0191_, w_1442_, w_2112_);
xor (w_0272_, new_in6[4], new_in18[4]);
nand (w_1473_, new_in4[4], w_1106_);
or (w_1271_, new_in21[3], w_2056_);
nand (w_2201_, w_1231_, w_0378_);
xor (w_0392_, new_in12[2], new_in15[0]);
nand (w_1799_, w_1398_, w_0250_);
xor (w_0962_, w_1989_, w_1342_);
xor (w_1950_, w_1571_, w_1737_);
nand (w_1108_, w_1131_, w_1832_);
nand (w_0280_, w_0263_, w_1468_);
xor (w_0093_, new_in7[2], new_in8[3]);
nand (w_0243_, new_in5[6], w_0053_);
and (w_0283_, new_in18[0], new_in20[1]);
or (w_1943_, new_in14[0], new_in22[1]);
nand (w_2010_, w_0345_, w_1462_);
nand (w_0931_, w_2061_, w_0894_);
or (w_1967_, w_1502_, w_2256_);
xor (w_0938_, w_1290_, w_1066_);
xor (w_0946_, w_0700_, w_1645_);
nand (w_0713_, w_0462_, w_1340_);
or (w_0483_, w_2093_, new_in1[0]);
xor (w_0514_, new_in20[6], w_1439_);
nor (new_out18[4], w_0170_, w_1229_);
xor (w_0811_, w_1744_, w_1128_);
or (w_0027_, w_1232_, w_2204_);
and (w_0829_, w_0098_, w_1749_);
nand (w_1237_, w_1520_, w_1735_);
nand (w_0142_, new_in1[4], new_in9[4]);
nand (w_1244_, new_in16[7], new_in22[0]);
and (w_1021_, new_in16[0], w_0244_);
xor (w_1034_, new_in19[4], new_in6[3]);
or (w_1251_, w_1627_, w_1300_);
nand (w_1483_, w_2270_, w_0217_);
nand (w_1639_, new_in16[7], w_0436_);
and (w_0460_, w_1473_, w_0076_);
nand (w_0558_, w_1839_, w_1920_);
nor (w_1603_, w_1231_, w_1952_);
nand (w_0637_, w_0757_, w_0545_);
nand (w_0375_, w_2106_, w_1081_);
and (w_2100_, new_in16[7], w_0154_);
xor (w_1674_, w_1091_, w_0592_);
xor (w_0436_, w_2288_, w_1125_);
or (w_0961_, w_2093_, w_2085_);
nand (w_1947_, new_in16[7], w_0784_);
or (w_1637_, w_2099_, w_2040_);
nand (w_1130_, new_in16[7], w_1089_);
not (w_2068_, new_in23[2]);
xor (w_1697_, new_in7[3], new_in15[3]);
xor (w_1463_, w_1479_, w_0580_);
nand (w_0521_, w_0700_, w_0423_);
xor (w_1595_, w_1752_, w_0743_);
nand (w_0270_, w_1847_, w_1612_);
xor (w_1984_, new_in20[3], w_0711_);
nand (w_1443_, w_1926_, w_0850_);
xor (w_0854_, w_0126_, w_1184_);
nand (w_1163_, w_2229_, w_0569_);
xor (w_1440_, w_1537_, w_0854_);
xor (w_0047_, new_in23[3], new_in6[3]);
nand (w_1436_, w_0368_, w_1936_);
xor (w_0855_, new_in22[3], new_in16[3]);
xor (w_2192_, new_in22[2], new_in16[2]);
nand (w_1044_, w_1231_, w_0021_);
xor (w_1201_, w_2313_, w_0149_);
xor (w_0895_, w_0351_, w_1910_);
and (w_0310_, w_0594_, w_0766_);
and (w_1722_, w_2098_, w_1344_);
nand (w_1500_, w_2184_, w_0657_);
xor (w_1747_, new_in22[0], new_in14[0]);
xor (w_1381_, new_in8[0], new_in1[0]);
xor (w_2240_, w_0489_, w_2303_);
xor (w_1017_, w_1791_, w_0051_);
nand (w_1318_, w_0882_, w_1257_);
nand (w_0728_, w_0263_, w_0510_);
nand (w_1932_, w_1231_, w_0952_);
nand (w_2059_, w_0136_, w_1482_);
nand (w_1400_, w_1231_, w_1870_);
xor (w_0059_, new_in4[3], new_in2[3]);
xor (w_1995_, new_in19[2], new_in17[2]);
nand (w_0327_, w_1465_, w_1682_);
nand (w_1306_, new_in20[5], w_1218_);
xor (w_0274_, w_2245_, w_1731_);
xor (w_1366_, w_0793_, w_0337_);
not (w_0458_, new_in16[0]);
or (w_1475_, w_0129_, w_0350_);
nand (w_0844_, w_1886_, w_0631_);
nand (w_0488_, w_1035_, w_1884_);
and (w_0162_, w_0649_, w_1309_);
and (new_out8[0], w_0438_, w_0109_);
nand (w_1102_, new_in5[6], w_0453_);
or (w_0447_, w_0144_, w_1891_);
xor (w_2253_, new_in7[5], new_in8[6]);
xor (w_0167_, w_2179_, w_0042_);
nand (w_1976_, new_in16[7], w_1074_);
nand (w_1838_, new_in10[8], w_0667_);
or (w_0442_, w_1231_, w_0773_);
xor (w_0443_, new_in23[4], new_in6[4]);
xor (w_0548_, w_0367_, w_2013_);
or (w_1514_, w_1052_, w_2226_);
nor (new_out14[2], w_1998_, w_1591_);
xor (w_1269_, w_0535_, w_1385_);
and (w_1520_, w_0741_, w_0090_);
or (w_1581_, w_0456_, w_1774_);
or (w_0341_, w_0759_, w_0068_);
or (w_1224_, w_0725_, w_0167_);
xor (w_0661_, new_in21[5], new_in3[5]);
nand (w_1902_, w_1234_, w_0611_);
xor (w_1934_, w_1247_, w_0207_);
nand (w_0984_, new_in21[1], new_in3[1]);
nor (w_1998_, w_1231_, w_0413_);
not (w_1663_, new_in1[2]);
nand (w_0857_, w_1234_, w_0477_);
and (w_1370_, new_in5[0], new_in9[1]);
xor (w_2194_, w_0652_, w_0196_);
xor (w_2256_, w_2175_, w_1097_);
xor (w_2015_, new_in21[3], new_in3[3]);
xor (w_0288_, w_2184_, w_1727_);
nand (w_1056_, w_1667_, w_0059_);
and (w_2109_, w_0281_, w_1122_);
or (w_0380_, w_2093_, w_1286_);
nand (w_0782_, w_1776_, w_0941_);
xor (w_0722_, w_0295_, w_0543_);
nand (w_1374_, w_2173_, w_2212_);
or (w_1382_, w_0920_, w_2032_);
xor (w_0549_, new_in14[2], new_in21[2]);
nand (w_1803_, new_in16[7], w_2073_);
nor (w_0796_, w_0793_, w_0337_);
not (w_1853_, w_1330_);
nand (w_0465_, w_1212_, w_1404_);
nand (w_0714_, new_in24[5], new_in2[5]);
nand (w_0219_, w_1937_, w_0180_);
nand (w_0018_, w_1873_, w_0320_);
and (new_out1[2], w_1101_, w_1223_);
xor (w_1621_, new_in14[2], new_in22[3]);
or (w_0827_, w_0263_, w_0445_);
or (w_1121_, w_1995_, w_0319_);
or (w_0639_, w_0212_, w_1589_);
xor (w_2172_, new_in1[2], new_in13[2]);
nand (w_0835_, w_0365_, w_2290_);
nand (w_0346_, w_2227_, w_2041_);
nand (w_0520_, w_0984_, w_0346_);
nand (w_0992_, new_in23[5], new_in6[5]);
xor (w_1207_, w_1532_, w_2224_);
nand (w_0266_, w_0880_, w_1656_);
and (w_0358_, new_in21[0], new_in20[1]);
nor (w_0837_, new_in13[3], w_2013_);
xor (w_0290_, new_in22[1], new_in16[1]);
and (w_1342_, new_in23[6], new_in12[6]);
xor (w_0139_, w_2130_, w_1901_);
xor (w_0994_, w_0608_, w_0301_);
xor (w_0873_, w_1485_, w_0179_);
xor (w_1831_, new_in4[0], new_in3[0]);
nor (w_0505_, w_0263_, w_1726_);
nand (w_0761_, w_0483_, w_1903_);
or (w_1188_, w_2057_, w_2208_);
xor (w_0244_, new_in3[0], w_0128_);
xor (w_1487_, new_in13[0], new_in13[1]);
nand (w_2116_, w_0499_, w_0665_);
or (w_1788_, w_1820_, w_2038_);
nand (w_0859_, w_0637_, w_2207_);
nand (w_1311_, w_1758_, w_0366_);
nand (w_1371_, w_0263_, w_1093_);
nand (new_out11[2], w_0273_, w_2002_);
and (w_0897_, w_0263_, w_0032_);
and (w_0113_, new_in5[6], w_1049_);
nand (w_1873_, w_1905_, w_0038_);
and (w_0510_, w_0442_, w_0463_);
xor (w_1135_, new_in6[6], new_in18[5]);
and (w_0212_, w_1928_, w_1156_);
nand (w_0774_, w_1231_, w_0716_);
and (w_1357_, w_1507_, w_0209_);
and (w_1180_, new_in7[0], new_in15[0]);
nand (w_1918_, w_1814_, w_2042_);
xor (w_0787_, new_in14[6], new_in21[6]);
nand (w_1380_, w_2136_, w_1009_);
and (w_1047_, w_0837_, w_1911_);
nand (w_1293_, w_0099_, w_0101_);
or (w_0132_, w_0729_, w_1280_);
nand (w_1290_, w_0987_, w_0731_);
xor (w_1307_, new_in19[3], new_in17[3]);
nand (w_0168_, w_0724_, w_1681_);
or (w_0418_, w_0283_, w_0822_);
xor (w_0145_, new_in1[5], new_in8[5]);
xor (w_1059_, w_0752_, w_1474_);
nand (w_0322_, w_1596_, w_1268_);
nand (w_0978_, w_1234_, w_2122_);
nand (w_0926_, w_1831_, w_0923_);
or (w_0013_, w_0255_, w_0033_);
nand (w_2270_, new_in20[3], w_0171_);
or (w_2202_, w_2255_, w_0305_);
nand (w_0349_, w_0331_, w_1391_);
xor (w_2076_, w_1226_, w_0392_);
nand (new_out12[5], w_1494_, w_0146_);
nand (w_1365_, w_0885_, w_0335_);
nand (w_0451_, new_in17[5], new_in10[5]);
not (w_0752_, new_in19[4]);
nand (w_1882_, new_in1[2], new_in8[1]);
nand (w_0009_, w_1234_, w_2091_);
nand (w_1147_, new_in5[6], w_1795_);
xor (w_0590_, w_0107_, w_0983_);
xor (w_2308_, w_0830_, w_1869_);
nand (w_1499_, w_0297_, w_1006_);
not (w_2026_, w_1538_);
nor (new_out18[5], w_2148_, w_1722_);
nand (w_1086_, w_1829_, w_0278_);
xor (w_1066_, new_in20[2], w_2138_);
xor (w_0289_, new_in19[3], new_in12[3]);
or (w_0815_, w_0429_, w_2231_);
and (new_out13[0], w_2267_, w_1688_);
xor (w_0792_, w_1566_, w_1909_);
xor (w_0775_, new_in18[2], new_in11[2]);
and (new_out11[4], w_2103_, w_1648_);
nand (w_1613_, w_0612_, w_0671_);
and (w_0539_, new_in20[0], w_2022_);
nand (w_1749_, w_1875_, w_1383_);
nand (w_2180_, w_0959_, w_2031_);
nand (w_1711_, w_1073_, w_0636_);
xor (w_0621_, w_1889_, w_1615_);
and (w_0295_, w_0768_, w_0527_);
nand (w_1824_, w_1313_, w_2269_);
nand (w_0967_, new_in16[2], w_1397_);
and (w_0061_, new_in5[6], w_0192_);
nand (w_1430_, w_0693_, w_1090_);
not (w_1338_, w_1508_);
and (w_2262_, w_1637_, w_1492_);
or (w_1437_, w_0263_, w_1366_);
nand (w_1255_, new_in3[2], w_1549_);
xor (w_0394_, w_1831_, w_2271_);
and (w_0014_, w_0923_, w_1514_);
nand (w_0750_, w_0215_, w_1263_);
xor (w_1656_, new_in20[5], w_1218_);
nand (new_out10[3], w_0034_, w_0924_);
xor (w_0126_, new_in19[4], new_in17[4]);
xor (w_1626_, w_1085_, w_0687_);
nand (w_2062_, w_1744_, w_1128_);
xor (w_1116_, new_in23[2], new_in12[2]);
nand (w_1640_, w_1312_, w_0293_);
nand (w_0254_, w_1231_, w_2107_);
and (w_0300_, new_in16[7], w_1730_);
nand (w_1228_, w_1681_, w_1182_);
nand (w_0339_, w_0263_, w_1392_);
nand (w_0189_, new_in22[1], new_in16[1]);
xor (w_0494_, w_1021_, w_0795_);
nand (w_0631_, w_1689_, w_0210_);
nand (w_0797_, w_0323_, w_0433_);
nand (w_2134_, new_in16[7], w_0002_);
xor (w_1721_, w_1414_, w_2321_);
nand (w_1786_, w_1502_, w_0237_);
xor (w_1693_, w_1352_, w_1605_);
or (w_1052_, w_1831_, w_2271_);
or (w_0841_, w_0680_, w_1559_);
nand (w_0830_, w_1575_, w_1541_);
nand (w_0748_, w_2193_, w_1215_);
nand (w_0814_, w_0432_, w_1561_);
nand (w_1112_, w_0712_, w_0977_);
nand (new_out11[3], w_2123_, w_1572_);
xor (w_1990_, new_in8[0], w_1705_);
nand (w_1134_, w_1628_, w_1816_);
and (w_1590_, w_1758_, w_1271_);
xor (w_2204_, w_1769_, w_0020_);
and (w_0049_, w_0110_, w_0933_);
or (w_0898_, new_in20[0], w_0422_);
xor (w_1850_, w_0667_, w_2078_);
xor (w_1496_, w_0215_, w_1840_);
nand (w_0552_, new_in16[7], w_1954_);
xor (w_0849_, w_1671_, w_1187_);
nand (w_0099_, w_0688_, w_2024_);
xor (w_1593_, new_in20[3], w_0171_);
nand (w_1706_, w_1205_, w_0512_);
and (w_0381_, new_in13[0], new_in24[0]);
nand (w_0430_, new_in21[3], new_in20[4]);
nand (w_1347_, new_in21[1], w_2001_);
nand (w_1782_, w_1588_, w_2189_);
nand (w_0553_, w_0142_, w_1935_);
or (w_1454_, w_0263_, w_1641_);
xor (w_1534_, new_in16[2], w_1202_);
nand (new_out16[5], w_0106_, w_0513_);
or (w_0467_, w_0574_, w_1584_);
and (w_1418_, w_0263_, w_2096_);
or (w_1523_, w_2323_, w_0016_);
or (w_0417_, w_0880_, w_1656_);
nand (w_0364_, w_0115_, w_1166_);
nand (w_2020_, w_1790_, w_1864_);
xor (w_0737_, w_1483_, w_2111_);
nand (new_out5[6], w_0927_, w_0554_);
xor (w_0401_, w_1587_, w_0185_);
xor (w_1262_, w_1455_, w_1301_);
nand (w_0389_, w_2093_, w_1957_);
nand (w_1826_, w_0131_, w_0420_);
xor (w_0355_, new_in1[3], w_1746_);
or (w_1813_, w_1752_, w_0743_);
nand (w_1189_, w_1725_, w_0762_);
xor (w_1295_, new_in9[2], new_in15[2]);
xor (w_1810_, w_1588_, w_2189_);
or (w_1929_, new_in20[0], w_2198_);
and (w_0609_, new_in23[4], new_in12[4]);
nand (w_0304_, w_0406_, w_1700_);
nand (w_1006_, w_1670_, w_0471_);
and (w_1930_, w_1631_, w_0057_);
xor (w_1845_, new_in17[0], new_in10[1]);
xor (w_2316_, w_0871_, w_0392_);
not (w_2210_, w_0215_);
nand (w_2044_, w_2191_, w_0964_);
xor (w_1774_, w_0423_, w_1019_);
or (w_1142_, w_1231_, w_1369_);
and (new_out17[5], w_1959_, w_0160_);
nand (w_0640_, w_1889_, w_0504_);
nand (w_1095_, w_0816_, w_0640_);
xor (w_1321_, w_0175_, w_1155_);
xor (w_0876_, w_1913_, w_0139_);
xor (w_1584_, new_in20[4], w_1781_);
xor (w_0262_, w_0376_, w_0881_);
xor (w_1871_, new_in14[5], new_in22[6]);
nand (w_0173_, w_0255_, w_0033_);
nand (w_0362_, w_1905_, w_2030_);
nand (w_1547_, w_2092_, w_0661_);
xor (w_0751_, w_1738_, w_1618_);
and (w_0077_, w_0263_, w_1102_);
and (w_0908_, w_0263_, w_2044_);
or (w_0846_, w_2124_, w_0155_);
nand (w_1388_, w_1443_, w_1411_);
xor (w_2226_, w_1499_, w_0684_);
xor (w_0179_, w_0374_, w_0755_);
nand (w_0643_, w_0357_, w_1616_);
xor (w_1913_, new_in19[0], new_in17[0]);
or (new_out5[0], w_2254_, w_1767_);
nand (w_0432_, w_1234_, w_2225_);
and (w_1470_, w_1052_, w_2226_);
nand (w_0331_, new_in17[1], new_in10[1]);
nand (w_1361_, w_0174_, w_1779_);
nand (new_out7[1], w_0776_, w_0875_);
nand (w_1184_, w_0216_, w_1001_);
or (w_0258_, w_0263_, w_2295_);
or (w_2250_, w_1171_, w_0197_);
xor (w_0511_, w_0118_, w_0060_);
or (w_1080_, w_2255_, w_1579_);
xor (w_2297_, new_in13[1], new_in24[1]);
nand (w_1692_, new_in16[7], w_1943_);
nand (w_1486_, w_1158_, w_1809_);
nand (w_0532_, w_1826_, w_1633_);
nand (w_0997_, w_1193_, w_1592_);
nand (w_1297_, w_1728_, w_2147_);
xor (w_0525_, w_1035_, w_1884_);
nand (w_0674_, w_0676_, w_1931_);
nand (w_0834_, new_in5[6], w_1460_);
and (w_1897_, w_0493_, w_1586_);
nand (w_1880_, w_1677_, w_0061_);
xor (w_0847_, w_1330_, w_1599_);
endmodule

module new_sub_module2(
    input wire new_in1,
    input wire new_in10,
    input wire new_in11,
    input wire new_in12,
    input wire new_in13,
    input wire new_in14,
    input wire new_in15,
    input wire new_in16,
    input wire new_in17,
    input wire new_in18,
    input wire new_in19,
    input wire new_in2,
    input wire new_in20,
    input wire new_in21,
    input wire new_in22,
    input wire new_in23,
    input wire new_in24,
    input wire new_in25,
    input wire new_in3,
    input wire new_in4,
    input wire new_in5,
    input wire new_in6,
    input wire new_in7,
    input wire new_in8,
    input wire new_in9,
    output wire new_out1,
    output wire new_out10,
    output wire new_out11,
    output wire new_out12,
    output wire new_out13,
    output wire new_out14,
    output wire new_out15,
    output wire new_out16,
    output wire new_out17,
    output wire new_out18,
    output wire new_out19,
    output wire new_out2,
    output wire new_out20,
    output wire new_out3,
    output wire new_out4,
    output wire new_out5,
    output wire new_out6,
    output wire new_out7,
    output wire new_out8,
    output wire new_out9
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
wire w_060_;
wire w_061_;
wire w_062_;
wire w_063_;
wire w_064_;
wire w_065_;
wire w_066_;
wire w_067_;
wire w_068_;
wire w_069_;
wire w_070_;
wire w_071_;
wire w_072_;
wire w_073_;
wire w_074_;
wire w_075_;
wire w_076_;
wire w_077_;
wire w_078_;
wire w_079_;
wire w_080_;
wire w_081_;
wire w_082_;
wire w_083_;
wire w_084_;
wire w_085_;
wire w_086_;
wire w_087_;
wire w_088_;
wire w_089_;
wire w_090_;
wire w_091_;
wire w_092_;
wire w_093_;
wire w_094_;
wire w_095_;
wire w_096_;
wire w_097_;
wire w_098_;
wire w_099_;
wire w_100_;
wire w_101_;
wire w_102_;
wire w_103_;
wire w_104_;
wire w_105_;
wire w_106_;
wire w_107_;
wire w_108_;
wire w_109_;
wire w_110_;
wire w_111_;
wire w_112_;
wire w_113_;
wire w_114_;
wire w_115_;
wire w_116_;
wire w_117_;
wire w_118_;
wire w_119_;
wire w_120_;
wire w_121_;
wire w_122_;
wire w_123_;
wire w_124_;
wire w_125_;
wire w_126_;
wire w_127_;
wire w_128_;
wire w_129_;
wire w_130_;
wire w_131_;
wire w_132_;
wire w_133_;
wire w_134_;
wire w_135_;
wire w_136_;
wire w_137_;
wire w_138_;
wire w_139_;
wire w_140_;
wire w_141_;
wire w_142_;
wire w_143_;
wire w_144_;
wire w_145_;
wire w_146_;
wire w_147_;
wire w_148_;
wire w_149_;
wire w_150_;
wire w_151_;
wire w_152_;
wire w_153_;
wire w_154_;
wire w_155_;
wire w_156_;
wire w_157_;
wire w_158_;
wire w_159_;
wire w_160_;
wire w_161_;
wire w_162_;
wire w_163_;
wire w_164_;
wire w_165_;
wire w_166_;
wire w_167_;
wire w_168_;
wire w_169_;
wire w_170_;
wire w_171_;
wire w_172_;
wire w_173_;
wire w_174_;
wire w_175_;
wire w_176_;
wire w_177_;
wire w_178_;
wire w_179_;
wire w_180_;
wire w_181_;
wire w_182_;
wire w_183_;
wire w_184_;
wire w_185_;
wire w_186_;
wire w_187_;
wire w_188_;
wire w_189_;
wire w_190_;
wire w_191_;
wire w_192_;
wire w_193_;
wire w_194_;
wire w_195_;
wire w_196_;
wire w_197_;
wire w_198_;
wire w_199_;
wire w_200_;
wire w_201_;
wire w_202_;
wire w_203_;
wire w_204_;
wire w_205_;
wire w_206_;
wire w_207_;
wire w_208_;
wire w_209_;
wire w_210_;
wire w_211_;
wire w_212_;
wire w_213_;
wire w_214_;
wire w_215_;
wire w_216_;
wire w_217_;
wire w_218_;
wire w_219_;
wire w_220_;
wire w_221_;
wire w_222_;
wire w_223_;
wire w_224_;
wire w_225_;
wire w_226_;
wire w_227_;
wire w_228_;
wire w_229_;
wire w_230_;
wire w_231_;
wire w_232_;
wire w_233_;
wire w_234_;
wire w_235_;
wire w_236_;
wire w_237_;
wire w_238_;
wire w_239_;
wire w_240_;
wire w_241_;
wire w_242_;
wire w_243_;
wire w_244_;
wire w_245_;
wire w_246_;
wire w_247_;
wire w_248_;
wire w_249_;
wire w_250_;
wire w_251_;
wire w_252_;
wire w_253_;
wire w_254_;
wire w_255_;
wire w_256_;
wire w_257_;
wire w_258_;
wire w_259_;
wire w_260_;
wire w_261_;
wire w_262_;
wire w_263_;
wire w_264_;
wire w_265_;
wire w_266_;
wire w_267_;
wire w_268_;
wire w_269_;
wire w_270_;
wire w_271_;
wire w_272_;
wire w_273_;
wire w_274_;
wire w_275_;
wire w_276_;
wire w_277_;
wire w_278_;
wire w_279_;
wire w_280_;
wire w_281_;
wire w_282_;
wire w_283_;
wire w_284_;
wire w_285_;
wire w_286_;
wire w_287_;
wire w_288_;
wire w_289_;
wire w_290_;
wire w_291_;
wire w_292_;
wire w_293_;
wire w_294_;
wire w_295_;
wire w_296_;
wire w_297_;
wire w_298_;
wire w_299_;
nor (w_072_, w_196_, w_000_);
nand (w_098_, w_199_, w_033_);
nand (w_082_, w_121_, w_291_);
and (w_003_, w_152_, w_128_);
and (w_047_, w_008_, w_052_);
nand (w_245_, w_196_, w_079_);
and (w_002_, w_054_, new_in9);
nor (w_235_, w_196_, w_102_);
nand (w_256_, w_161_, w_017_);
nand (w_094_, w_157_, w_076_);
nand (w_004_, w_227_, w_011_);
nand (w_241_, w_196_, w_122_);
or (w_069_, w_227_, w_011_);
xor (w_266_, w_029_, w_179_);
nand (w_195_, w_143_, w_124_);
and (w_176_, new_in12, new_in6);
xor (w_196_, new_in8, new_in4);
and (w_240_, w_244_, w_227_);
nand (w_130_, w_143_, w_146_);
or (w_055_, w_196_, w_111_);
nand (new_out1, w_042_, w_057_);
nand (new_out9, w_180_, w_110_);
nand (new_out7, w_212_, w_153_);
nor (w_217_, w_029_, w_179_);
nand (w_023_, w_200_, w_064_);
nand (w_254_, w_200_, w_094_);
not (w_054_, new_in8);
nand (w_071_, w_119_, w_275_);
xor (w_171_, w_142_, w_011_);
nand (w_095_, w_157_, w_261_);
and (w_085_, w_111_, w_244_);
nand (w_158_, w_121_, w_113_);
nand (w_115_, w_027_, w_121_);
or (w_211_, w_121_, w_060_);
nor (w_001_, w_094_, w_261_);
nand (w_060_, w_200_, w_091_);
and (w_253_, w_143_, w_181_);
and (w_272_, w_142_, w_037_);
or (w_205_, w_064_, w_089_);
nand (w_163_, w_004_, w_162_);
nand (w_099_, w_143_, w_259_);
nand (w_284_, w_142_, w_200_);
nand (w_057_, w_199_, w_243_);
nand (w_182_, w_088_, w_240_);
and (w_150_, w_296_, w_025_);
or (w_073_, w_027_, w_000_);
and (w_262_, w_199_, w_142_);
nand (w_090_, w_064_, w_014_);
and (w_200_, new_in4, w_189_);
nand (w_108_, w_266_, w_244_);
nand (w_120_, w_229_, w_129_);
xor (w_076_, new_in19, new_in22);
and (w_079_, w_111_, w_064_);
and (w_169_, new_in3, w_141_);
nand (new_out13, w_050_, w_276_);
nand (w_238_, w_121_, w_190_);
nand (w_114_, w_043_, w_091_);
xor (w_012_, w_029_, w_157_);
nand (w_128_, w_266_, w_091_);
nand (w_214_, w_027_, w_075_);
nand (w_101_, w_199_, w_094_);
xor (w_215_, w_043_, w_142_);
xor (w_165_, w_227_, w_157_);
not (w_221_, new_in13);
and (new_out6, w_021_, w_026_);
nand (w_151_, w_199_, w_092_);
nand (w_203_, w_090_, w_250_);
and (w_246_, w_115_, w_209_);
nand (w_089_, w_196_, w_167_);
xor (w_164_, w_200_, w_091_);
xor (w_207_, w_227_, w_027_);
nand (w_007_, w_027_, w_200_);
nand (new_out12, w_074_, w_270_);
and (w_144_, w_223_, w_290_);
nand (w_287_, w_199_, w_298_);
and (w_132_, new_in14, new_in5);
and (w_077_, w_121_, w_089_);
and (w_064_, w_297_, new_in24);
and (w_059_, w_143_, w_194_);
or (w_040_, w_004_, w_060_);
and (w_044_, w_029_, w_121_);
nand (w_194_, w_004_, w_060_);
nand (w_154_, w_196_, w_280_);
nand (w_018_, w_213_, w_255_);
or (w_223_, w_196_, w_288_);
nand (w_188_, w_232_, w_154_);
and (w_258_, w_220_, w_036_);
and (w_159_, w_199_, w_055_);
and (w_278_, w_214_, w_202_);
and (w_075_, w_244_, w_070_);
nand (w_153_, w_143_, w_147_);
nand (w_056_, w_244_, w_171_);
nand (w_066_, w_027_, w_279_);
nand (w_065_, w_121_, w_015_);
or (w_232_, w_196_, w_246_);
and (w_091_, w_157_, w_076_);
nand (w_027_, w_134_, w_248_);
nor (w_237_, w_196_, w_044_);
nand (new_out19, w_192_, w_178_);
nand (w_127_, w_121_, w_018_);
and (w_045_, w_043_, w_011_);
or (w_010_, w_196_, w_136_);
nand (w_134_, new_in8, w_111_);
nand (w_036_, w_244_, w_046_);
nand (w_062_, w_222_, w_069_);
nand (w_078_, w_143_, w_164_);
xor (w_219_, w_298_, w_020_);
nand (w_000_, w_297_, new_in24);
and (w_020_, w_227_, w_142_);
nand (w_177_, w_199_, w_112_);
nand (w_019_, w_200_, w_011_);
or (w_186_, w_200_, w_187_);
nand (w_005_, w_196_, w_019_);
or (w_139_, w_196_, w_106_);
nand (w_290_, w_196_, w_060_);
nand (w_138_, w_199_, w_048_);
nand (w_048_, w_234_, w_245_);
and (w_265_, w_196_, w_043_);
and (w_141_, new_in25, new_in18);
nand (w_247_, w_196_, w_251_);
and (w_277_, w_289_, w_148_);
nand (w_061_, w_227_, w_200_);
nand (new_out3, w_024_, w_295_);
or (w_096_, w_029_, w_115_);
nand (w_192_, w_199_, w_030_);
nand (w_183_, w_121_, w_091_);
nand (w_295_, w_199_, w_144_);
or (w_022_, w_227_, w_091_);
nand (w_122_, w_254_, w_053_);
and (w_043_, new_in10, new_in16);
nand (w_049_, w_143_, w_219_);
nand (new_out16, w_197_, w_010_);
and (w_160_, w_266_, w_011_);
and (w_226_, w_233_, w_177_);
xor (w_014_, w_027_, w_170_);
and (w_136_, w_098_, w_252_);
and (w_068_, w_103_, w_239_);
or (w_034_, w_196_, w_150_);
and (w_105_, w_244_, w_022_);
nand (w_216_, w_196_, w_062_);
or (w_280_, w_157_, w_087_);
nand (w_093_, w_261_, w_107_);
nand (w_097_, w_142_, w_000_);
or (w_263_, w_157_, w_176_);
or (w_250_, w_014_, w_061_);
nand (w_028_, w_142_, w_085_);
or (w_296_, w_043_, w_108_);
nand (new_out15, w_117_, w_099_);
nand (w_166_, w_157_, w_236_);
nand (w_107_, w_027_, w_157_);
xor (w_111_, w_043_, w_179_);
nand (w_152_, w_142_, w_094_);
nand (w_104_, w_064_, w_125_);
xor (w_267_, w_142_, w_064_);
nand (w_233_, w_244_, w_273_);
nand (w_123_, w_249_, w_101_);
nand (w_197_, w_196_, w_269_);
nand (w_086_, w_116_, w_095_);
xor (w_201_, w_266_, w_014_);
nand (w_210_, w_121_, w_277_);
or (w_230_, w_196_, w_047_);
or (w_281_, w_196_, w_109_);
nand (w_255_, w_014_, w_292_);
nand (w_270_, w_199_, w_188_);
nand (w_024_, w_244_, w_263_);
and (new_out11, w_274_, w_005_);
nor (w_102_, w_134_, w_142_);
or (w_016_, w_001_, w_236_);
nand (w_252_, w_244_, w_084_);
or (w_174_, w_196_, w_126_);
nand (new_out20, w_210_, w_051_);
nand (new_out14, w_006_, w_158_);
and (w_162_, w_196_, w_298_);
nand (w_110_, w_143_, w_294_);
nand (w_243_, w_038_, w_238_);
and (w_179_, new_in11, new_in20);
nand (w_030_, w_230_, w_241_);
nor (w_035_, w_227_, w_287_);
nand (w_190_, w_293_, w_083_);
and (w_084_, w_027_, w_170_);
nand (new_out17, w_108_, w_149_);
nand (new_out4, w_138_, w_056_);
nand (w_257_, w_040_, w_059_);
nand (new_out5, w_155_, w_082_);
nand (w_083_, w_027_, w_072_);
nand (w_191_, w_143_, w_242_);
and (w_067_, w_078_, w_100_);
nand (w_206_, w_027_, w_215_);
nand (w_239_, w_121_, w_012_);
nand (w_299_, w_196_, w_203_);
and (w_063_, w_197_, w_031_);
nand (w_117_, w_121_, w_071_);
nand (w_038_, w_143_, w_041_);
or (w_119_, w_196_, w_286_);
nand (w_220_, w_043_, w_199_);
nand (w_092_, w_266_, w_094_);
or (w_218_, w_227_, w_064_);
and (w_009_, w_127_, w_049_);
nand (w_053_, w_091_, w_264_);
xor (w_142_, w_132_, w_184_);
nand (w_231_, w_121_, w_079_);
nand (w_146_, w_081_, w_224_);
nand (w_155_, w_143_, w_271_);
nor (w_032_, w_279_, w_035_);
xor (w_261_, w_064_, w_014_);
nand (w_109_, w_168_, w_285_);
xor (w_133_, w_142_, w_091_);
nand (w_170_, new_in12, new_in6);
nand (w_222_, w_227_, w_000_);
and (new_out2, w_195_, w_039_);
xor (w_271_, w_027_, w_091_);
and (w_031_, w_199_, w_135_);
nand (w_167_, w_142_, w_157_);
nand (w_131_, w_121_, w_123_);
nand (w_224_, w_043_, w_227_);
and (w_236_, w_064_, w_094_);
nand (w_148_, w_196_, w_114_);
xor (w_070_, w_043_, w_091_);
and (w_185_, w_094_, w_014_);
nand (w_006_, w_143_, w_201_);
nand (w_285_, w_143_, w_206_);
and (w_173_, w_043_, w_157_);
or (w_234_, w_196_, w_067_);
nand (w_249_, w_244_, w_086_);
or (w_051_, w_121_, w_137_);
and (w_292_, w_029_, w_244_);
nand (w_276_, w_131_, w_283_);
nand (w_161_, w_211_, w_237_);
xor (w_172_, w_227_, w_045_);
or (w_113_, w_105_, w_063_);
nand (w_124_, w_167_, w_116_);
nand (w_129_, w_199_, w_068_);
or (w_274_, w_196_, w_120_);
nand (w_242_, w_097_, w_104_);
nand (w_259_, w_282_, w_228_);
or (w_260_, w_196_, w_226_);
nand (w_106_, w_257_, w_096_);
or (w_046_, w_142_, w_058_);
nand (w_178_, w_244_, w_118_);
nand (w_199_, new_in17, new_in6);
nand (w_149_, w_139_, w_013_);
and (w_126_, w_140_, w_065_);
nand (w_015_, w_151_, w_066_);
xor (w_189_, new_in7, new_in1);
xor (w_294_, w_023_, w_185_);
nand (new_out10, w_174_, w_193_);
nand (w_187_, new_in17, w_147_);
nand (w_100_, w_227_, w_121_);
or (w_225_, w_196_, w_258_);
nand (w_042_, w_244_, w_198_);
nand (w_298_, new_in4, w_189_);
nand (w_074_, w_105_, w_268_);
nand (w_282_, w_111_, w_298_);
nand (w_033_, w_191_, w_183_);
nand (w_157_, w_156_, w_187_);
and (w_279_, w_244_, w_261_);
nand (w_145_, w_247_, w_260_);
nand (w_029_, new_in10, new_in16);
nand (w_135_, w_073_, w_235_);
nand (w_248_, w_142_, w_002_);
nand (w_268_, w_227_, w_091_);
or (w_289_, w_196_, w_032_);
xor (w_011_, w_027_, w_176_);
and (w_264_, w_142_, w_064_);
nand (w_052_, w_143_, w_172_);
nand (w_181_, w_007_, w_272_);
xor (w_118_, w_111_, w_027_);
or (w_026_, w_196_, w_009_);
or (w_041_, w_079_, w_160_);
and (w_143_, new_in24, new_in3);
and (w_184_, w_221_, new_in2);
nand (w_039_, w_121_, w_278_);
nand (w_212_, w_034_, w_077_);
nand (w_198_, w_186_, w_061_);
not (w_297_, new_in23);
nand (new_out18, w_175_, w_281_);
nand (w_208_, w_019_, w_282_);
nand (w_112_, w_266_, w_014_);
xor (w_269_, w_298_, w_173_);
nand (w_175_, w_196_, w_016_);
nand (w_121_, new_in24, new_in3);
and (w_017_, w_199_, w_216_);
and (w_204_, new_in21, new_in15);
nand (w_291_, w_299_, w_225_);
xor (w_273_, w_217_, w_027_);
or (w_213_, w_244_, w_118_);
nand (w_229_, w_244_, w_218_);
or (w_116_, w_064_, w_157_);
nand (w_202_, w_163_, w_159_);
or (w_228_, w_227_, w_298_);
nand (w_168_, w_182_, w_080_);
xor (w_147_, w_200_, w_064_);
nand (w_275_, w_196_, w_093_);
or (w_088_, w_111_, w_157_);
nand (w_021_, w_196_, w_166_);
or (w_140_, w_121_, w_284_);
and (w_080_, w_121_, w_287_);
xor (w_251_, w_157_, w_020_);
nor (w_283_, w_196_, w_253_);
nand (w_293_, w_133_, w_265_);
or (w_156_, new_in17, w_284_);
nand (w_180_, w_121_, w_145_);
nand (w_081_, w_029_, w_267_);
nand (new_out8, w_028_, w_256_);
or (w_125_, w_111_, w_227_);
nand (w_193_, w_196_, w_165_);
nor (w_286_, w_075_, w_262_);
nand (w_050_, w_196_, w_125_);
xor (w_058_, w_111_, w_157_);
and (w_013_, w_199_, w_205_);
nand (w_008_, w_121_, w_157_);
and (w_227_, w_204_, w_169_);
or (w_037_, w_027_, w_200_);
and (w_087_, w_043_, w_142_);
nand (w_209_, w_143_, w_208_);
nand (w_288_, w_130_, w_231_);
or (w_025_, w_244_, w_207_);
nand (w_103_, w_143_, w_003_);
and (w_244_, new_in17, new_in6);
xor (w_137_, w_142_, w_107_);
endmodule

module new_sub_module3(
    input wire [1:0] new_in1,
    input wire [1:0] new_in10,
    input wire [1:0] new_in11,
    input wire [1:0] new_in12,
    input wire [1:0] new_in13,
    input wire [1:0] new_in14,
    input wire [1:0] new_in15,
    input wire [1:0] new_in16,
    input wire [1:0] new_in17,
    input wire [1:0] new_in18,
    input wire [1:0] new_in19,
    input wire [1:0] new_in2,
    input wire [1:0] new_in20,
    input wire [1:0] new_in3,
    input wire [1:0] new_in4,
    input wire [1:0] new_in5,
    input wire [1:0] new_in6,
    input wire [1:0] new_in7,
    input wire [1:0] new_in8,
    input wire [1:0] new_in9,
    output wire [3:0] new_out1,
    output wire [3:0] new_out10,
    output wire [3:0] new_out11,
    output wire [3:0] new_out12,
    output wire [3:0] new_out13,
    output wire [3:0] new_out14,
    output wire [3:0] new_out15,
    output wire [3:0] new_out2,
    output wire [3:0] new_out3,
    output wire [3:0] new_out4,
    output wire [3:0] new_out5,
    output wire [3:0] new_out6,
    output wire [3:0] new_out7,
    output wire [3:0] new_out8,
    output wire [3:0] new_out9
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
nand (w_0284_, w_0185_, w_0512_);
nand (w_0404_, w_0858_, w_0282_);
or (w_0559_, w_0220_, w_0823_);
xor (w_0645_, w_0644_, w_0362_);
xor (w_0308_, new_in10[1], new_in12[1]);
xor (w_0537_, w_0611_, w_0519_);
xor (w_0503_, w_0357_, w_0687_);
xor (w_0074_, new_in19[0], new_in12[0]);
xor (w_0027_, w_0386_, w_0259_);
nand (w_0688_, w_0824_, w_0570_);
or (w_0780_, w_0824_, w_0159_);
nand (w_0606_, w_0695_, w_0649_);
nand (w_0504_, new_in11[1], w_0694_);
xor (w_0699_, w_0581_, w_0460_);
nand (w_0928_, w_0908_, w_0040_);
nand (w_0480_, new_in11[1], w_0377_);
nand (w_0215_, w_0186_, w_0738_);
and (w_0834_, w_0220_, w_0695_);
nand (w_0565_, w_0336_, w_0925_);
nand (new_out10[0], w_0363_, w_0544_);
and (w_0133_, w_0665_, w_0773_);
and (new_out11[0], w_0333_, w_0598_);
nand (w_0109_, w_0841_, w_0099_);
xor (w_0165_, w_0880_, w_0699_);
nand (w_0188_, w_0220_, w_0241_);
xor (w_0194_, new_in20[0], new_in19[0]);
nand (w_0226_, new_in13[1], w_0220_);
nand (w_0409_, w_0614_, w_0561_);
not (w_0600_, w_0525_);
nand (w_0575_, w_0297_, w_0441_);
xor (w_0660_, new_in11[1], new_in2[1]);
nand (w_0231_, w_0758_, w_0647_);
xor (w_0232_, new_in11[1], w_0623_);
xor (w_0923_, w_0298_, w_0376_);
and (w_0420_, new_in16[0], w_0665_);
or (w_0751_, w_0336_, w_0172_);
nand (w_0296_, w_0756_, w_0506_);
nand (w_0513_, w_0023_, w_0244_);
nand (w_0450_, w_0701_, w_0696_);
xor (w_0472_, w_0939_, w_0017_);
xor (w_0806_, w_0788_, w_0921_);
nand (new_out6[3], w_0774_, w_0310_);
xor (w_0056_, w_0279_, w_0604_);
nand (w_0359_, w_0834_, w_0399_);
xor (w_0269_, w_0464_, w_0577_);
nand (w_0690_, w_0679_, w_0876_);
xor (w_0901_, new_in4[1], new_in2[0]);
nand (w_0185_, new_in11[1], w_0623_);
and (w_0052_, new_in11[1], new_in8[1]);
nand (w_0616_, w_0008_, w_0105_);
nand (w_0933_, new_in11[0], new_in2[0]);
nand (w_0558_, w_0181_, w_0199_);
or (w_0845_, w_0824_, w_0198_);
nand (w_0440_, w_0008_, w_0289_);
nand (w_0327_, new_in20[0], new_in2[1]);
xor (w_0649_, w_0541_, w_0723_);
nand (w_0557_, w_0775_, w_0583_);
xor (w_0366_, new_in11[1], new_in4[1]);
xor (w_0490_, w_0109_, w_0640_);
xor (w_0137_, w_0124_, w_0916_);
or (w_0184_, w_0349_, w_0339_);
xor (w_0196_, new_in1[0], new_in13[0]);
and (w_0449_, w_0285_, w_0671_);
and (new_out3[3], w_0035_, w_0475_);
nand (w_0003_, w_0824_, w_0019_);
nand (w_0096_, w_0599_, new_in18[0]);
nand (w_0453_, w_0273_, w_0669_);
xor (w_0481_, new_in20[1], w_0550_);
nand (w_0841_, new_in1[1], new_in17[1]);
xor (w_0677_, w_0700_, w_0507_);
nand (w_0434_, w_0336_, w_0909_);
xor (w_0103_, w_0514_, w_0421_);
xor (w_0740_, w_0279_, new_in15[0]);
and (w_0224_, new_in4[0], new_in17[0]);
xor (w_0238_, w_0420_, w_0848_);
xor (w_0678_, w_0567_, w_0787_);
nand (w_0819_, w_0514_, w_0421_);
or (w_0140_, w_0336_, w_0367_);
nand (w_0605_, w_0613_, w_0207_);
or (w_0412_, w_0336_, w_0622_);
and (w_0516_, new_in11[0], new_in17[0]);
and (new_out2[1], w_0295_, w_0136_);
or (w_0000_, w_0352_, w_0829_);
nand (w_0119_, new_in7[1], new_in18[1]);
nand (w_0750_, w_0341_, w_0088_);
and (w_0797_, w_0725_, w_0068_);
nand (w_0361_, w_0692_, w_0132_);
nand (w_0601_, w_0043_, w_0702_);
and (w_0346_, w_0243_, w_0128_);
nand (w_0917_, w_0003_, w_0249_);
nand (w_0680_, w_0824_, w_0453_);
nand (w_0873_, w_0305_, w_0240_);
nand (w_0093_, w_0212_, w_0084_);
nand (w_0799_, w_0892_, w_0157_);
nand (w_0893_, w_0060_, w_0413_);
xor (w_0778_, new_in10[1], new_in14[1]);
or (w_0043_, w_0336_, w_0027_);
nand (w_0181_, new_in17[1], new_in8[1]);
and (w_0255_, w_0852_, new_in9[1]);
xor (w_0146_, w_0218_, w_0918_);
nand (w_0692_, new_in10[1], w_0833_);
xor (w_0805_, w_0650_, w_0285_);
nand (w_0010_, w_0858_, w_0742_);
or (w_0728_, w_0824_, w_0553_);
nand (w_0505_, w_0686_, w_0568_);
nand (w_0837_, w_0695_, w_0543_);
and (w_0072_, w_0220_, w_0564_);
nand (w_0081_, w_0516_, w_0535_);
nand (w_0104_, w_0841_, w_0341_);
and (w_0831_, new_in6[0], w_0220_);
nand (w_0217_, w_0008_, w_0778_);
nand (w_0256_, w_0685_, w_0660_);
nand (w_0863_, w_0824_, w_0818_);
nand (w_0240_, w_0336_, w_0798_);
nand (new_out4[1], w_0881_, w_0034_);
and (new_out15[2], w_0276_, w_0272_);
and (w_0506_, w_0336_, w_0674_);
nand (w_0907_, w_0195_, w_0415_);
nand (w_0903_, w_0090_, w_0476_);
and (w_0551_, w_0485_, w_0446_);
xor (w_0426_, new_in18[0], new_in12[0]);
xor (w_0339_, new_in10[1], new_in17[1]);
nand (w_0365_, w_0695_, w_0390_);
xor (w_0595_, w_0231_, w_0180_);
nor (w_0005_, w_0008_, w_0336_);
xor (w_0916_, w_0762_, w_0174_);
nand (w_0161_, new_in6[0], new_in7[0]);
nand (w_0919_, w_0336_, w_0393_);
or (w_0488_, w_0153_, w_0579_);
nand (w_0493_, w_0365_, w_0389_);
nand (w_0158_, w_0769_, w_0754_);
nand (new_out1[3], w_0190_, w_0451_);
nand (w_0311_, w_0695_, w_0872_);
or (w_0410_, w_0744_, w_0755_);
and (new_out6[2], w_0839_, w_0615_);
xor (w_0499_, w_0650_, w_0019_);
and (w_0549_, new_in3[0], w_0592_);
nand (w_0617_, w_0631_, w_0352_);
nand (w_0760_, w_0042_, w_0382_);
and (w_0867_, new_in1[0], new_in2[0]);
nand (w_0437_, w_0824_, w_0878_);
nand (w_0850_, w_0824_, w_0794_);
or (w_0588_, w_0336_, w_0855_);
nand (w_0247_, w_0505_, w_0525_);
and (w_0292_, w_0858_, w_0854_);
nand (w_0111_, new_in8[0], w_0858_);
xor (w_0904_, w_0775_, w_0766_);
or (w_0943_, w_0220_, w_0901_);
or (w_0735_, w_0609_, w_0805_);
xor (w_0457_, w_0285_, w_0671_);
nand (w_0594_, new_in7[0], new_in18[0]);
nand (w_0145_, w_0858_, w_0757_);
or (w_0885_, new_in10[1], w_0833_);
nand (w_0141_, w_0097_, w_0518_);
nand (w_0211_, w_0336_, w_0361_);
xor (w_0847_, new_in4[0], w_0345_);
or (w_0358_, w_0582_, w_0094_);
or (w_0839_, w_0220_, w_0682_);
xor (w_0198_, new_in10[0], new_in14[0]);
nand (w_0920_, w_0905_, w_0009_);
nand (w_0044_, w_0735_, w_0533_);
xor (w_0535_, new_in11[1], new_in17[1]);
nand (w_0243_, w_0221_, w_0255_);
nand (w_0064_, w_0858_, w_0143_);
nand (w_0079_, w_0430_, w_0341_);
nand (w_0489_, w_0025_, w_0092_);
xor (w_0854_, new_in10[1], new_in20[1]);
xor (w_0176_, new_in10[0], new_in20[0]);
or (w_0566_, w_0578_, w_0705_);
or (w_0273_, w_0695_, w_0150_);
nand (w_0338_, w_0211_, w_0348_);
nand (w_0474_, new_in6[0], new_in10[0]);
nand (w_0817_, w_0925_, w_0797_);
not (w_0613_, new_in18[1]);
nand (w_0173_, w_0394_, w_0827_);
nand (w_0078_, w_0824_, w_0448_);
nand (w_0897_, w_0299_, w_0321_);
nand (w_0814_, w_0858_, w_0840_);
nor (w_0125_, w_0876_, w_0555_);
nand (w_0560_, w_0824_, w_0830_);
or (w_0200_, new_in1[1], new_in13[1]);
nand (w_0421_, w_0342_, w_0069_);
nand (w_0286_, w_0216_, w_0246_);
xor (w_0514_, new_in6[0], new_in20[0]);
xor (w_0041_, w_0619_, w_0727_);
nand (w_0717_, w_0386_, w_0259_);
or (w_0021_, w_0220_, w_0406_);
xor (w_0223_, w_0462_, w_0325_);
nand (w_0482_, w_0695_, w_0698_);
xor (w_0828_, w_0737_, w_0820_);
xor (w_0679_, w_0867_, w_0710_);
or (w_0126_, w_0791_, w_0842_);
nand (w_0784_, w_0484_, w_0617_);
xor (w_0880_, w_0665_, w_0773_);
or (w_0563_, w_0449_, w_0672_);
xor (w_0843_, w_0485_, w_0392_);
xor (w_0647_, w_0775_, w_0876_);
nand (w_0403_, w_0434_, w_0596_);
nand (new_out11[2], w_0811_, w_0652_);
nand (w_0343_, w_0813_, w_0699_);
or (w_0118_, new_in11[0], new_in2[0]);
xor (w_0413_, w_0536_, w_0913_);
or (w_0393_, w_0220_, w_0183_);
nand (w_0135_, w_0858_, w_0056_);
nand (w_0374_, w_0939_, w_0017_);
xor (w_0895_, w_0285_, w_0019_);
nand (w_0869_, w_0188_, w_0064_);
or (w_0114_, new_in10[1], w_0008_);
nand (w_0369_, w_0695_, w_0074_);
nand (w_0618_, w_0314_, w_0171_);
nand (w_0057_, w_0343_, w_0897_);
nand (w_0193_, w_0008_, w_0937_);
nand (w_0794_, w_0638_, w_0919_);
nand (w_0351_, w_0637_, w_0277_);
xor (w_0935_, w_0194_, w_0082_);
or (w_0695_, new_in16[0], new_in5[1]);
xor (w_0473_, new_in5[1], w_0200_);
and (w_0567_, new_in1[0], new_in11[0]);
xor (w_0675_, w_0002_, w_0048_);
nand (new_out1[2], w_0175_, w_0139_);
nand (w_0058_, w_0729_, w_0127_);
nand (w_0556_, w_0718_, w_0569_);
nand (w_0719_, w_0153_, w_0579_);
nand (new_out8[1], w_0708_, w_0066_);
xor (w_0331_, new_in11[0], new_in13[0]);
nand (w_0621_, w_0586_, new_in12[0]);
nand (w_0761_, w_0459_, w_0317_);
xor (w_0370_, w_0061_, w_0497_);
and (w_0389_, w_0824_, w_0771_);
nand (w_0030_, w_0494_, w_0747_);
xor (w_0712_, new_in6[1], w_0483_);
nand (w_0648_, w_0858_, w_0375_);
nand (w_0414_, w_0341_, w_0806_);
nand (w_0628_, w_0274_, w_0815_);
xor (w_0597_, new_in1[0], new_in17[0]);
nand (w_0399_, new_in18[0], w_0392_);
and (w_0639_, w_0658_, w_0235_);
nand (w_0192_, w_0304_, w_0030_);
nand (w_0724_, w_0858_, w_0234_);
nand (w_0151_, w_0858_, w_0260_);
nand (new_out14[1], w_0222_, w_0584_);
or (w_0295_, w_0220_, w_0435_);
not (w_0871_, w_0325_);
nand (w_0236_, w_0220_, w_0498_);
nand (new_out1[0], w_0691_, w_0385_);
nor (w_0233_, w_0695_, w_0936_);
nand (w_0899_, w_0573_, w_0184_);
nand (w_0632_, w_0008_, w_0334_);
nand (w_0737_, w_0474_, w_0374_);
not (w_0510_, new_in8[0]);
and (w_0921_, w_0841_, w_0161_);
nand (w_0199_, w_0037_, w_0110_);
nand (w_0280_, w_0858_, w_0862_);
xor (w_0773_, new_in11[1], new_in8[1]);
xor (w_0641_, new_in20[1], w_0178_);
nand (w_0883_, new_in20[0], new_in19[0]);
nand (w_0020_, w_0858_, w_0103_);
and (w_0028_, w_0857_, w_0071_);
or (w_0857_, w_0336_, w_0935_);
and (w_0380_, new_in7[0], w_0220_);
or (w_0008_, w_0255_, w_0694_);
or (w_0328_, w_0336_, w_0783_);
and (w_0936_, new_in6[1], w_0220_);
and (new_out7[1], w_0853_, w_0890_);
or (w_0025_, w_0824_, w_0481_);
or (w_0046_, w_0824_, w_0462_);
and (w_0589_, w_0786_, w_0247_);
or (w_0376_, w_0775_, w_0766_);
and (w_0536_, w_0524_, w_0566_);
nand (w_0772_, w_0163_, w_0087_);
nand (w_0065_, w_0325_, w_0392_);
xor (w_0466_, new_in6[0], new_in19[0]);
xor (w_0143_, new_in8[1], w_0678_);
and (new_out2[0], w_0162_, w_0941_);
nand (w_0716_, w_0695_, w_0522_);
nand (w_0075_, w_0695_, w_0400_);
or (w_0468_, new_in20[1], w_0695_);
nand (w_0139_, w_0336_, w_0799_);
nand (w_0353_, w_0115_, w_0165_);
and (w_0268_, w_0824_, w_0425_);
or (w_0447_, w_0336_, w_0091_);
nand (w_0801_, new_in10[0], w_0745_);
or (w_0401_, w_0336_, w_0418_);
and (w_0439_, w_0220_, w_0739_);
xor (w_0024_, new_in17[1], w_0462_);
nand (w_0568_, w_0558_, w_0636_);
nand (w_0701_, w_0298_, w_0131_);
nand (w_0433_, w_0336_, w_0672_);
nand (w_0864_, w_0414_, w_0770_);
xor (w_0525_, new_in6[1], new_in12[1]);
or (w_0718_, w_0220_, w_0387_);
nand (w_0138_, w_0117_, w_0574_);
xor (w_0397_, new_in6[1], new_in18[1]);
and (w_0900_, new_in1[1], w_0220_);
nand (w_0865_, w_0220_, w_0469_);
nand (w_0324_, w_0336_, w_0107_);
xor (w_0120_, new_in9[0], w_0736_);
xor (w_0400_, new_in4[1], w_0219_);
nand (w_0478_, w_0824_, w_0173_);
nand (w_0070_, w_0824_, w_0051_);
nand (w_0379_, w_0336_, w_0016_);
nand (w_0492_, w_0515_, w_0072_);
and (w_0768_, w_0050_, w_0528_);
xor (w_0775_, w_0465_, w_0318_);
or (w_0049_, w_0163_, w_0087_);
or (w_0562_, new_in1[0], new_in2[0]);
nand (w_0896_, w_0220_, w_0626_);
nand (w_0381_, w_0662_, w_0779_);
or (w_0555_, w_0650_, w_0019_);
xor (w_0271_, new_in3[0], w_0592_);
nand (w_0838_, w_0220_, w_0542_);
or (w_0208_, w_0336_, w_0350_);
nand (w_0195_, w_0008_, w_0270_);
nand (w_0225_, w_0167_, w_0417_);
or (w_0937_, new_in7[0], new_in18[0]);
or (w_0001_, w_0805_, w_0503_);
nand (w_0190_, w_0336_, w_0039_);
nand (w_0942_, w_0858_, w_0611_);
nand (w_0249_, w_0008_, w_0116_);
nand (w_0098_, w_0634_, w_0759_);
xor (w_0318_, new_in10[0], new_in12[0]);
xor (w_0159_, w_0115_, w_0165_);
or (w_0669_, w_0336_, w_0677_);
xor (w_0861_, w_0681_, w_0191_);
nand (w_0889_, w_0332_, new_in2[1]);
nand (w_0812_, w_0341_, w_0329_);
xor (w_0091_, new_in13[1], new_in17[1]);
xor (w_0477_, new_in6[1], w_0610_);
xor (w_0875_, w_0174_, w_0261_);
nand (w_0715_, new_in12[1], w_0292_);
nand (w_0347_, w_0581_, w_0460_);
xor (w_0915_, w_0868_, w_0527_);
xor (w_0171_, new_in9[1], w_0460_);
xor (w_0152_, new_in13[0], new_in17[0]);
xor (w_0387_, w_0758_, w_0647_);
nor (w_0859_, new_in7[1], new_in19[1]);
or (w_0424_, w_0824_, w_0683_);
nand (w_0932_, w_0432_, w_0242_);
xor (w_0511_, w_0462_, w_0392_);
or (w_0691_, w_0336_, w_0152_);
nand (w_0117_, w_0187_, w_0373_);
or (w_0105_, new_in7[1], new_in18[1]);
nand (w_0136_, w_0220_, w_0287_);
nand (w_0908_, w_0442_, w_0291_);
and (w_0178_, w_0319_, w_0452_);
nand (new_out14[0], w_0471_, w_0910_);
xor (w_0055_, w_0511_, w_0517_);
nand (w_0796_, w_0336_, w_0360_);
nand (w_0790_, w_0858_, w_0120_);
xor (w_0213_, new_in3[0], w_0703_);
and (w_0294_, w_0220_, w_0489_);
nand (new_out10[3], w_0364_, w_0763_);
and (new_out5[2], w_0149_, w_0303_);
and (w_0519_, w_0344_, w_0819_);
or (w_0090_, w_0695_, w_0012_);
nand (w_0252_, w_0858_, w_0137_);
nand (new_out8[3], w_0673_, w_0616_);
or (w_0573_, new_in10[1], w_0332_);
nand (w_0730_, new_in1[1], new_in11[1]);
nand (w_0039_, w_0018_, w_0715_);
not (w_0168_, w_0186_);
xor (w_0543_, new_in13[1], new_in8[1]);
nand (w_0931_, w_0008_, w_0562_);
xor (w_0309_, w_0325_, w_0668_);
nor (w_0452_, new_in4[0], new_in4[1]);
nand (w_0471_, w_0220_, w_0932_);
nand (w_0486_, w_0220_, w_0849_);
xor (w_0019_, w_0037_, w_0110_);
and (w_0128_, w_0220_, w_0504_);
xor (w_0636_, new_in6[0], new_in12[0]);
nand (w_0248_, new_in20[1], new_in19[1]);
nand (w_0348_, w_0695_, w_0590_);
nand (w_0892_, new_in12[0], w_0229_);
nand (w_0383_, w_0679_, w_0699_);
nand (w_0187_, w_0488_, w_0866_);
nand (w_0402_, w_0858_, w_0275_);
nand (w_0655_, new_in18[1], w_0834_);
xor (w_0650_, new_in17[0], new_in8[0]);
nand (w_0122_, w_0411_, w_0502_);
not (w_0745_, new_in19[0]);
xor (w_0418_, new_in9[0], w_0671_);
or (w_0638_, w_0336_, w_0331_);
nand (w_0642_, w_0695_, w_0602_);
xor (w_0687_, w_0019_, w_0679_);
nand (w_0846_, w_0332_, w_0462_);
xor (w_0592_, new_in11[0], new_in8[0]);
or (w_0175_, w_0336_, w_0466_);
xor (w_0390_, w_0325_, w_0125_);
nand (w_0396_, w_0326_, w_0102_);
or (w_0707_, w_0220_, w_0861_);
and (w_0578_, w_0279_, new_in13[0]);
nand (w_0250_, new_in11[1], new_in2[1]);
nand (w_0112_, w_0045_, w_0914_);
nand (w_0659_, w_0824_, w_0874_);
and (w_0608_, w_0336_, w_0726_);
nand (w_0704_, w_0552_, w_0302_);
xor (w_0191_, new_in18[1], w_0207_);
xor (w_0077_, new_in20[0], new_in2[0]);
nor (w_0654_, w_0879_, w_0251_);
and (w_0386_, w_0285_, w_0019_);
nand (w_0038_, w_0852_, w_0699_);
nand (w_0333_, w_0695_, w_0802_);
and (w_0320_, w_0858_, w_0106_);
nand (w_0378_, w_0824_, w_0900_);
and (w_0088_, new_in17[0], w_0592_);
nand (w_0419_, w_0824_, w_0189_);
or (w_0076_, w_0597_, w_0362_);
nand (w_0603_, w_0898_, w_0268_);
nand (w_0063_, w_0699_, w_0630_);
and (w_0630_, new_in2[1], w_0834_);
nor (w_0336_, new_in16[0], new_in5[1]);
nand (w_0827_, w_0858_, w_0828_);
xor (w_0781_, w_0019_, w_0431_);
and (w_0502_, w_0008_, w_0013_);
nand (w_0033_, w_0803_, w_0169_);
xor (w_0587_, w_0592_, w_0671_);
and (w_0722_, new_in8[1], w_0858_);
nand (w_0739_, w_0695_, w_0194_);
nor (w_0886_, new_in1[0], new_in13[0]);
nand (w_0022_, new_in9[1], w_0460_);
xor (w_0714_, w_0879_, w_0251_);
xor (w_0727_, new_in18[1], new_in10[1]);
and (w_0619_, w_0350_, w_0141_);
or (w_0007_, w_0336_, w_0895_);
nand (new_out3[2], w_0205_, w_0020_);
nand (w_0911_, new_in16[1], w_0052_);
and (w_0277_, w_0220_, w_0680_);
nand (w_0107_, w_0812_, w_0943_);
nand (w_0572_, w_0194_, w_0082_);
nand (w_0475_, w_0493_, w_0004_);
or (w_0124_, w_0664_, w_0490_);
nand (w_0313_, w_0635_, w_0194_);
and (w_0314_, new_in9[0], w_0671_);
xor (w_0377_, w_0880_, w_0019_);
and (w_0405_, w_0118_, w_0927_);
or (w_0720_, w_0824_, w_0355_);
nand (new_out4[2], w_0863_, w_0257_);
and (w_0368_, w_0220_, w_0046_);
nand (w_0517_, w_0383_, w_0258_);
nand (new_out11[3], w_0307_, w_0075_);
xor (w_0611_, new_in6[1], new_in20[1]);
xor (w_0422_, w_0477_, w_0155_);
nor (w_0816_, w_0220_, w_0196_);
nand (new_out4[0], w_0227_, w_0427_);
xor (w_0862_, w_0631_, w_0352_);
nand (w_0532_, w_0220_, w_0059_);
nand (w_0276_, w_0220_, w_0443_);
nand (w_0534_, w_0462_, w_0871_);
and (w_0218_, w_0810_, w_0121_);
and (w_0287_, w_0210_, w_0632_);
and (w_0684_, w_0419_, w_0580_);
nand (w_0212_, w_0912_, w_0011_);
nand (w_0815_, w_0695_, w_0844_);
and (w_0037_, new_in17[0], new_in8[0]);
xor (w_0802_, w_0745_, w_0699_);
or (w_0461_, w_0261_, w_0033_);
nand (new_out5[0], w_0444_, w_0532_);
xor (w_0264_, w_0060_, w_0413_);
nand (w_0807_, w_0824_, w_0876_);
nand (new_out1[1], w_0209_, w_0447_);
nand (w_0265_, w_0858_, w_0213_);
nand (w_0626_, w_0704_, w_0311_);
or (w_0142_, w_0336_, w_0509_);
nand (w_0067_, w_0109_, w_0640_);
nand (w_0538_, w_0624_, w_0540_);
xor (w_0267_, w_0654_, w_0031_);
nand (w_0051_, w_0627_, w_0944_);
nand (new_out3[0], w_0724_, w_0547_);
nand (w_0470_, w_0557_, w_0316_);
xor (w_0703_, new_in17[0], new_in2[0]);
xor (w_0260_, w_0397_, w_0633_);
and (w_0445_, w_0585_, w_0096_);
nand (w_0709_, w_0465_, w_0318_);
nand (w_0006_, w_0079_, w_0340_);
nand (w_0627_, w_0858_, w_0753_);
nand (w_0609_, w_0220_, w_0008_);
and (w_0809_, w_0083_, w_0378_);
nand (w_0767_, w_0646_, w_0468_);
nand (w_0127_, w_0366_, w_0722_);
not (w_0813_, w_0876_);
or (w_0524_, w_0221_, new_in13[1]);
nand (w_0756_, w_0858_, w_0714_);
and (w_0229_, w_0858_, w_0176_);
or (w_0726_, w_0609_, w_0663_);
nand (w_0326_, w_0824_, w_0767_);
xor (w_0392_, w_0635_, w_0194_);
or (w_0272_, w_0220_, w_0835_);
nand (w_0515_, w_0336_, w_0429_);
nor (w_0824_, w_0255_, w_0694_);
xor (w_0713_, w_0381_, w_0230_);
xor (w_0012_, w_0352_, w_0829_);
nand (w_0144_, new_in13[0], new_in8[0]);
or (w_0465_, w_0052_, w_0133_);
and (w_0395_, w_0670_, w_0408_);
and (w_0822_, w_0248_, w_0738_);
or (w_0624_, w_0925_, w_0797_);
nand (w_0774_, w_0220_, w_0575_);
xor (w_0234_, new_in8[0], w_0840_);
and (new_out12[0], w_0501_, w_0751_);
and (w_0009_, w_0119_, w_0105_);
or (w_0239_, w_0220_, w_0438_);
and (w_0204_, w_0220_, w_0424_);
xor (w_0657_, w_0599_, w_0899_);
nand (w_0580_, w_0008_, w_0523_);
and (new_out6[0], w_0135_, w_0492_);
xor (w_0527_, new_in10[1], new_in19[1]);
nand (w_0777_, w_0625_, w_0928_);
and (w_0721_, w_0341_, w_0479_);
xor (w_0682_, w_0284_, w_0653_);
and (w_0810_, w_0781_, w_0301_);
nand (new_out13[0], w_0796_, w_0856_);
or (w_0798_, w_0220_, w_0055_);
nor (w_0851_, w_0312_, w_0679_);
nand (w_0528_, w_0325_, w_0005_);
and (w_0693_, new_in18[1], new_in10[1]);
and (w_0153_, new_in15[0], w_0431_);
nand (w_0702_, w_0336_, w_0639_);
and (w_0102_, w_0220_, w_0217_);
xor (w_0116_, new_in15[0], w_0671_);
xor (w_0509_, w_0775_, w_0392_);
xor (w_0150_, w_0202_, w_0643_);
xor (w_0629_, w_0349_, w_0339_);
and (w_0665_, new_in11[0], new_in8[0]);
nand (w_0026_, w_0008_, w_0740_);
nand (w_0016_, w_0860_, w_0782_);
or (w_0197_, w_0336_, w_0587_);
nand (w_0156_, w_0001_, w_0891_);
xor (w_0345_, w_0168_, w_0822_);
nand (w_0877_, w_0336_, w_0760_);
xor (w_0698_, new_in17[0], w_0679_);
xor (w_0508_, new_in1[0], w_0592_);
nand (w_0771_, w_0336_, w_0041_);
xor (w_0134_, w_0668_, w_0589_);
nand (w_0749_, w_0929_, w_0800_);
and (w_0084_, w_0594_, w_0937_);
xor (w_0237_, new_in8[1], w_0281_);
nand (w_0130_, w_0645_, w_0803_);
and (w_0497_, w_0732_, w_0593_);
and (new_out11[1], w_0140_, w_0324_);
and (w_0388_, w_0695_, w_0772_);
nand (w_0095_, w_0695_, w_0734_);
nand (w_0487_, w_0026_, w_0437_);
nand (w_0101_, w_0300_, w_0330_);
and (new_out7[0], w_0006_, w_0197_);
not (w_0262_, new_in16[1]);
nand (w_0830_, w_0486_, w_0145_);
nand (w_0706_, w_0804_, w_0353_);
and (w_0054_, w_0695_, w_0089_);
and (w_0288_, w_0220_, w_0283_);
or (w_0415_, w_0008_, w_0589_);
xor (w_0017_, new_in6[0], new_in10[0]);
xor (w_0522_, new_in10[0], new_in17[0]);
nand (w_0906_, w_0410_, w_0320_);
or (w_0856_, w_0336_, w_0933_);
nand (w_0335_, new_in1[0], w_0824_);
xor (w_0040_, w_0876_, w_0462_);
xor (w_0048_, new_in18[0], new_in20[1]);
not (w_0384_, w_0668_);
nand (w_0108_, w_0008_, w_0370_);
xor (w_0671_, new_in4[0], new_in13[0]);
xor (w_0330_, new_in20[0], new_in2[1]);
xor (w_0855_, w_0298_, w_0345_);
nand (w_0770_, w_0858_, w_0269_);
xor (w_0742_, w_0733_, w_0859_);
nand (new_out8[2], w_0193_, w_0731_);
and (w_0485_, w_0038_, w_0488_);
nand (w_0205_, w_0323_, w_0204_);
nand (w_0069_, w_0224_, w_0406_);
nand (w_0547_, w_0938_, w_0894_);
xor (w_0281_, w_0224_, w_0406_);
xor (w_0753_, new_in7[0], w_0047_);
nand (w_0129_, new_in6[0], new_in18[0]);
nand (w_0429_, w_0008_, w_0597_);
xor (w_0844_, w_0876_, w_0555_);
nand (w_0725_, w_0462_, w_0392_);
nand (w_0372_, w_0906_, w_0608_);
nand (w_0501_, w_0336_, w_0809_);
xor (w_0087_, new_in6[0], w_0668_);
xor (w_0325_, w_0505_, w_0600_);
xor (w_0653_, w_0192_, w_0426_);
nand (w_0241_, w_0924_, w_0433_);
nand (w_0708_, w_0824_, w_0338_);
nand (w_0316_, w_0101_, w_0832_);
nand (w_0697_, w_0791_, w_0842_);
and (new_out5[1], w_0707_, w_0170_);
xor (w_0306_, w_0279_, new_in4[0]);
nand (w_0625_, w_0876_, w_0462_);
xor (w_0876_, w_0558_, w_0636_);
nand (w_0853_, w_0032_, w_0293_);
nand (w_0696_, w_0858_, w_0675_);
and (new_out6[1], w_0559_, w_0423_);
nand (w_0416_, new_in11[1], new_in17[1]);
nand (w_0789_, w_0546_, w_0233_);
or (w_0425_, new_in4[1], w_0695_);
xor (w_0925_, w_0384_, w_0345_);
xor (w_0523_, new_in14[0], w_0285_);
or (w_0154_, w_0676_, w_0223_);
xor (w_0764_, w_0345_, w_0589_);
nand (w_0651_, w_0695_, w_0693_);
nand (w_0582_, new_in11[0], w_0312_);
xor (w_0147_, w_0612_, w_0713_);
and (w_0341_, w_0220_, w_0008_);
and (w_0349_, new_in10[0], w_0312_);
xor (w_0495_, new_in18[0], w_0597_);
and (w_0293_, w_0336_, w_0104_);
xor (w_0602_, w_0893_, w_0915_);
xor (w_0747_, new_in8[1], new_in2[1]);
nand (w_0930_, w_0412_, w_0789_);
and (w_0430_, new_in1[0], new_in17[0]);
nand (w_0633_, w_0129_, w_0148_);
and (w_0529_, w_0858_, w_0697_);
or (w_0940_, new_in10[0], w_0008_);
nand (w_0662_, new_in18[0], new_in12[0]);
and (w_0732_, new_in13[1], new_in8[1]);
nand (w_0686_, new_in6[0], new_in12[0]);
nand (w_0222_, w_0780_, w_0166_);
xor (w_0577_, new_in5[1], new_in12[1]);
and (w_0866_, w_0008_, w_0719_);
nand (w_0228_, w_0336_, w_0864_);
nand (w_0591_, w_0008_, w_0904_);
or (w_0938_, w_0419_, w_0405_);
xor (w_0463_, new_in1[1], new_in13[1]);
nand (w_0808_, w_0220_, w_0286_);
nand (w_0073_, w_0008_, w_0146_);
and (w_0744_, w_0689_, w_0126_);
and (w_0540_, w_0858_, w_0817_);
nand (w_0310_, w_0858_, w_0147_);
xor (w_0672_, w_0679_, w_0699_);
nand (w_0254_, w_0336_, w_0538_);
and (new_out7[2], w_0372_, w_0142_);
nand (w_0743_, w_0336_, w_0761_);
nand (w_0018_, w_0220_, w_0122_);
xor (w_0230_, w_0613_, new_in12[1]);
nand (w_0929_, w_0049_, w_0388_);
xor (w_0842_, new_in16[1], new_in8[1]);
nand (w_0571_, w_0858_, w_0508_);
nand (w_0752_, new_in4[0], w_0858_);
nand (w_0484_, new_in17[1], new_in2[1]);
nand (w_0769_, new_in7[0], new_in10[0]);
and (w_0059_, w_0884_, w_0007_);
nor (w_0723_, w_0700_, w_0507_);
not (w_0644_, w_0597_);
xor (w_0438_, w_0409_, w_0775_);
nand (w_0407_, w_0008_, w_0781_);
xor (w_0251_, new_in7[0], new_in19[0]);
nand (w_0610_, w_0119_, w_0920_);
xor (w_0462_, w_0212_, w_0084_);
xor (w_0836_, w_0314_, w_0171_);
nand (w_0763_, w_0008_, w_0923_);
xor (w_0352_, new_in17[1], new_in2[1]);
nand (w_0209_, w_0336_, w_0058_);
nand (w_0323_, w_0824_, w_0628_);
nand (w_0042_, w_0858_, w_0514_);
nand (w_0354_, w_0065_, w_0576_);
nand (w_0596_, w_0695_, w_0422_);
and (w_0620_, new_in11[0], w_0604_);
xor (w_0180_, w_0298_, w_0325_);
nand (w_0821_, new_in18[0], w_0008_);
xor (w_0334_, new_in14[1], w_0679_);
nand (new_out12[2], w_0369_, w_0556_);
nand (w_0612_, w_0284_, w_0653_);
nand (w_0615_, w_0461_, w_0439_);
nand (new_out14[2], w_0351_, w_0790_);
or (w_0160_, w_0336_, w_0250_);
nand (w_0912_, new_in1[1], new_in2[1]);
nand (w_0253_, w_0942_, w_0888_);
or (w_0661_, w_0851_, w_0024_);
or (w_0189_, w_0336_, w_0650_);
xor (w_0666_, w_0810_, w_0121_);
xor (w_0848_, new_in16[1], w_0052_);
nand (w_0849_, w_0398_, w_0565_);
xor (w_0668_, w_0905_, w_0009_);
nand (w_0123_, w_0220_, w_0917_);
or (w_0729_, w_0609_, w_0036_);
or (w_0902_, w_0695_, w_0703_);
xor (w_0840_, new_in4[0], new_in17[0]);
nand (w_0498_, w_0659_, w_0440_);
nand (w_0924_, w_0695_, w_0629_);
nand (w_0307_, w_0336_, w_0450_);
nand (w_0833_, w_0258_, w_0563_);
not (w_0586_, new_in5[0]);
nand (w_0157_, w_0156_, w_0721_);
nand (w_0011_, w_0867_, w_0710_);
nand (new_out13[3], w_0651_, w_0086_);
and (w_0300_, new_in4[1], new_in2[0]);
nand (w_0305_, w_0695_, w_0264_);
nand (w_0363_, w_0824_, w_0776_);
nand (w_0491_, w_0220_, w_0487_);
xor (w_0174_, new_in6[1], new_in7[1]);
and (w_0163_, w_0846_, w_0661_);
xor (w_0623_, w_0494_, w_0747_);
or (w_0544_, w_0592_, w_0824_);
nand (w_0939_, w_0416_, w_0081_);
or (w_0275_, w_0196_, w_0463_);
xor (w_0455_, new_in2[1], w_0113_);
nand (new_out2[3], w_0648_, w_0467_);
nand (w_0576_, w_0057_, w_0062_);
nand (w_0329_, new_in17[1], w_0880_);
or (w_0169_, w_0640_, w_0076_);
nand (w_0552_, w_0008_, w_0455_);
nand (w_0758_, w_0480_, w_0358_);
and (w_0803_, w_0008_, w_0336_);
xor (w_0539_, new_in6[1], new_in19[1]);
or (w_0394_, w_0345_, w_0655_);
nand (w_0459_, w_0220_, w_0513_);
xor (w_0085_, w_0777_, w_0309_);
nand (new_out14[3], w_0236_, w_0010_);
nand (w_0106_, w_0744_, w_0755_);
nand (w_0441_, w_0803_, w_0875_);
nand (w_0099_, w_0430_, w_0362_);
xor (w_0734_, new_in19[1], new_in12[1]);
xor (w_0029_, w_0445_, w_0397_);
xor (w_0362_, new_in1[1], new_in17[1]);
nand (w_0244_, new_in18[1], w_0008_);
xor (w_0062_, w_0325_, w_0392_);
nand (w_0910_, w_0858_, w_0711_);
nand (w_0035_, w_0858_, w_0537_);
or (w_0428_, w_0336_, w_0807_);
and (w_0541_, new_in10[1], new_in12[1]);
nand (w_0782_, w_0824_, w_0380_);
xor (w_0047_, new_in11[0], new_in17[0]);
nand (w_0786_, new_in6[1], new_in12[1]);
and (new_out10[1], w_0053_, w_0728_);
xor (w_0622_, w_0851_, w_0024_);
and (w_0004_, w_0220_, w_0108_);
nand (w_0561_, w_0549_, w_0667_);
and (w_0593_, new_in19[0], new_in12[0]);
and (w_0469_, w_0821_, w_0335_);
nand (w_0245_, w_0700_, w_0709_);
nand (w_0652_, w_0336_, w_0470_);
nand (new_out15[0], w_0265_, w_0491_);
nand (w_0360_, w_0123_, w_0814_);
nand (w_0258_, w_0449_, w_0672_);
xor (w_0823_, w_0620_, w_0232_);
or (w_0427_, new_in4[0], w_0824_);
nand (w_0342_, new_in4[1], new_in17[1]);
nand (w_0884_, w_0336_, w_0112_);
nand (w_0170_, w_0220_, w_0601_);
or (w_0014_, w_0536_, w_0913_);
not (w_0548_, w_0057_);
nand (w_0089_, w_0676_, w_0223_);
and (w_0373_, w_0220_, w_0807_);
or (w_0546_, w_0879_, w_0402_);
nand (w_0186_, w_0883_, w_0313_);
or (w_0274_, w_0695_, w_0203_);
or (w_0898_, w_0336_, w_0836_);
nand (w_0656_, w_0008_, w_0843_);
and (w_0278_, w_0328_, w_0902_);
nand (w_0317_, w_0858_, w_0595_);
nand (w_0201_, w_0008_, w_0144_);
nand (w_0283_, w_0695_, w_0460_);
and (w_0357_, w_0650_, w_0285_);
or (w_0411_, w_0156_, w_0085_);
nand (w_0776_, w_0530_, w_0482_);
nand (w_0530_, w_0336_, w_0015_);
and (w_0762_, w_0161_, w_0067_);
not (w_0599_, new_in6[0]);
xor (w_0757_, new_in12[1], w_0765_);
nand (w_0673_, w_0824_, w_0870_);
xor (w_0711_, w_0586_, w_0886_);
and (w_0894_, w_0220_, w_0201_);
and (w_0436_, w_0336_, w_0752_);
and (w_0115_, w_0592_, w_0671_);
nand (w_0301_, w_0897_, w_0793_);
nand (w_0826_, w_0824_, w_0903_);
nand (w_0689_, w_0262_, new_in8[1]);
nand (w_0080_, w_0567_, w_0787_);
and (new_out9[2], w_0688_, w_0266_);
nand (w_0795_, w_0428_, w_0368_);
xor (w_0663_, w_0841_, w_0161_);
not (w_0446_, w_0392_);
not (w_0279_, new_in11[0]);
and (new_out2[2], w_0239_, w_0795_);
nand (w_0032_, w_0126_, w_0529_);
xor (w_0683_, w_0732_, w_0593_);
and (w_0261_, w_0640_, w_0076_);
not (w_0685_, w_0933_);
xor (w_0207_, w_0430_, w_0362_);
nor (w_0829_, w_0312_, new_in2[0]);
nand (new_out13[1], w_0160_, w_0138_);
xor (w_0285_, new_in1[0], new_in2[0]);
nand (new_out9[1], w_0078_, w_0720_);
and (w_0060_, w_0331_, w_0882_);
xor (w_0640_, new_in6[0], new_in7[0]);
nand (w_0888_, w_0220_, w_0907_);
nand (w_0214_, w_0336_, w_0457_);
xor (w_0913_, new_in10[0], new_in19[0]);
nand (w_0266_, w_0008_, w_0666_);
or (w_0736_, new_in7[0], new_in19[0]);
xor (w_0182_, w_0822_, w_0572_);
and (w_0550_, new_in20[0], new_in2[0]);
nand (w_0382_, w_0220_, w_0741_);
nand (w_0607_, w_0420_, w_0848_);
nand (w_0423_, w_0130_, w_0288_);
nand (w_0408_, w_0706_, w_0509_);
xor (w_0321_, w_0813_, w_0699_);
or (w_0890_, w_0336_, w_0165_);
and (w_0569_, w_0336_, w_0865_);
nand (new_out8[0], w_0850_, w_0931_);
nand (w_0741_, w_0656_, w_0164_);
or (w_0914_, new_in11[0], w_0008_);
nand (w_0785_, new_in13[1], new_in4[1]);
xor (w_0202_, new_in6[0], new_in18[0]);
not (w_0319_, new_in20[0]);
nand (w_0257_, w_0008_, w_0922_);
xor (w_0667_, new_in3[1], w_0880_);
or (w_0533_, w_0111_, w_0306_);
nand (w_0385_, w_0336_, w_0044_);
nand (w_0350_, new_in18[0], new_in10[0]);
and (w_0464_, w_0621_, w_0410_);
nand (w_0868_, w_0801_, w_0014_);
not (w_0332_, new_in17[1]);
nand (w_0263_, w_0858_, w_0267_);
xor (w_0121_, w_0548_, w_0062_);
or (w_0637_, w_0824_, w_0746_);
xor (w_0110_, new_in17[1], new_in8[1]);
nand (w_0909_, w_0226_, w_0263_);
or (w_0793_, w_0299_, w_0321_);
xor (w_0934_, w_0933_, w_0660_);
nand (w_0874_, w_0206_, w_0606_);
xor (w_0036_, w_0805_, w_0503_);
xor (w_0435_, w_0549_, w_0667_);
xor (w_0765_, w_0158_, w_0500_);
xor (w_0100_, w_0516_, w_0535_);
and (w_0443_, w_0496_, w_0845_);
nand (w_0216_, w_0695_, w_0657_);
xor (w_0882_, w_0578_, w_0705_);
and (w_0507_, w_0911_, w_0607_);
xor (w_0456_, new_in7[0], new_in10[0]);
and (new_out10[2], w_0591_, w_0749_);
xor (w_0375_, w_0322_, w_0298_);
nand (new_out7[3], w_0228_, w_0588_);
nand (w_0635_, w_0785_, w_0347_);
xor (w_0579_, new_in15[1], w_0699_);
or (w_0476_, w_0336_, w_0238_);
nand (w_0113_, new_in20[1], w_0550_);
and (w_0927_, w_0336_, w_0933_);
and (w_0061_, new_in19[1], new_in12[1]);
xor (w_0031_, new_in7[1], new_in19[1]);
xor (w_0460_, new_in13[1], new_in4[1]);
or (w_0585_, w_0202_, w_0643_);
nand (w_0634_, w_0336_, w_0934_);
and (w_0858_, new_in3[1], new_in14[0]);
or (w_0164_, w_0008_, w_0325_);
not (w_0312_, new_in17[0]);
xor (w_0553_, w_0592_, w_0880_);
or (w_0034_, w_0824_, w_0454_);
xor (w_0872_, w_0371_, w_0134_);
nand (w_0881_, w_0824_, w_0869_);
nand (new_out5[3], w_0896_, w_0252_);
xor (w_0748_, w_0582_, w_0094_);
or (w_0658_, w_0221_, w_0008_);
and (w_0766_, w_0592_, w_0880_);
nand (w_0520_, w_0571_, w_0838_);
nand (w_0219_, w_0248_, w_0215_);
or (w_0451_, w_0336_, w_0539_);
nand (w_0297_, w_0695_, w_0822_);
xor (w_0820_, new_in6[1], new_in10[1]);
and (new_out15[1], w_0280_, w_0315_);
nand (w_0598_, w_0750_, w_0436_);
and (w_0132_, w_0858_, w_0885_);
xor (w_0454_, new_in4[0], new_in4[1]);
xor (w_0891_, w_0908_, w_0040_);
and (w_0155_, w_0554_, w_0049_);
xor (w_0458_, w_0664_, w_0490_);
nand (w_0315_, w_0603_, w_0346_);
and (w_0092_, w_0336_, w_0940_);
nand (w_0731_, w_0824_, w_0873_);
nand (w_0646_, w_0695_, w_0182_);
and (w_0832_, w_0858_, w_0179_);
nand (w_0531_, w_0154_, w_0054_);
nand (w_0083_, new_in17[0], w_0858_);
nand (new_out12[3], w_0743_, w_0095_);
nand (w_0442_, w_0019_, w_0679_);
nand (new_out13[2], w_0208_, w_0877_);
xor (w_0355_, w_0781_, w_0301_);
and (w_0494_, new_in8[0], new_in2[0]);
nand (w_0584_, w_0858_, w_0473_);
xor (w_0918_, w_0354_, w_0764_);
xor (w_0590_, w_0331_, w_0882_);
and (w_0681_, new_in18[0], w_0644_);
or (w_0391_, new_in4[0], w_0695_);
or (w_0926_, w_0220_, w_0472_);
and (w_0800_, w_0824_, w_0296_);
and (w_0694_, new_in15[1], w_0733_);
nand (new_out4[3], w_0560_, w_0177_);
or (w_0738_, new_in20[1], new_in19[1]);
or (w_0356_, new_in1[1], new_in2[1]);
and (w_0631_, new_in17[0], new_in2[0]);
and (w_0791_, new_in16[0], w_0510_);
or (w_0674_, new_in13[0], w_0858_);
and (w_0340_, w_0336_, w_0111_);
xor (w_0282_, new_in7[1], w_0100_);
nand (w_0818_, w_0808_, w_0337_);
nand (w_0700_, new_in10[0], new_in12[0]);
and (w_0302_, w_0336_, w_0114_);
nand (w_0779_, w_0192_, w_0426_);
nand (w_0788_, new_in6[1], new_in7[1]);
xor (w_0787_, new_in1[1], new_in11[1]);
xor (w_0203_, w_0097_, w_0518_);
xor (w_0094_, w_0221_, w_0377_);
or (w_0479_, w_0001_, w_0891_);
nand (new_out9[3], w_0478_, w_0073_);
and (w_0581_, new_in4[0], new_in13[0]);
xor (w_0710_, new_in1[1], new_in2[1]);
nand (w_0149_, w_0858_, w_0458_);
nand (w_0303_, w_0531_, w_0294_);
nand (w_0299_, w_0019_, w_0431_);
and (w_0574_, w_0336_, w_0021_);
xor (w_0755_, new_in5[0], new_in12[0]);
nand (w_0227_, w_0824_, w_0520_);
nand (w_0496_, w_0824_, w_0028_);
or (w_0015_, w_0831_, w_0816_);
or (w_0811_, w_0336_, w_0847_);
nand (w_0002_, w_0327_, w_0101_);
not (w_0733_, new_in9[1]);
nand (w_0432_, w_0824_, w_0278_);
nand (new_out3[1], w_0225_, w_0521_);
nand (w_0053_, w_0824_, w_0930_);
nand (w_0148_, w_0202_, w_0784_);
nand (w_0905_, w_0594_, w_0093_);
not (w_0221_, new_in11[1]);
nand (w_0941_, w_0220_, w_0684_);
or (w_0177_, w_0824_, w_0641_);
or (w_0526_, w_0681_, w_0191_);
nand (w_0564_, w_0695_, w_0671_);
nand (w_0290_, new_in2[0], w_0220_);
xor (w_0298_, w_0245_, w_0308_);
xor (w_0545_, w_0887_, w_0456_);
and (w_0676_, w_0690_, w_0717_);
xor (w_0259_, w_0679_, w_0876_);
xor (w_0172_, new_in13[0], new_in8[0]);
and (w_0417_, w_0220_, w_0792_);
nand (w_0614_, new_in3[1], w_0880_);
xor (w_0705_, new_in11[1], new_in13[1]);
nand (w_0887_, w_0730_, w_0080_);
nand (w_0097_, w_0250_, w_0256_);
nand (w_0344_, new_in6[0], new_in20[0]);
xor (w_0183_, new_in10[0], w_0457_);
nand (w_0235_, w_0008_, w_0077_);
nand (w_0068_, w_0511_, w_0517_);
xor (w_0270_, w_0551_, w_0345_);
nand (w_0570_, w_0926_, w_0359_);
xor (w_0500_, new_in7[1], new_in10[1]);
or (w_0050_, w_0824_, w_0668_);
or (w_0179_, w_0300_, w_0330_);
nand (w_0246_, w_0336_, w_0511_);
xor (w_0783_, new_in16[0], w_0665_);
nand (w_0554_, w_0599_, w_0668_);
and (w_0583_, w_0008_, w_0831_);
xor (w_0406_, new_in4[1], new_in17[1]);
and (w_0643_, w_0000_, w_0889_);
nand (w_0664_, w_0605_, w_0526_);
xor (w_0604_, new_in8[0], new_in2[0]);
nand (new_out9[0], w_0070_, w_0407_);
xor (w_0289_, w_0395_, w_0855_);
not (w_0431_, w_0671_);
or (w_0210_, w_0336_, w_0003_);
nand (new_out12[1], w_0837_, w_0379_);
nand (w_0220_, new_in3[1], new_in14[0]);
xor (w_0825_, new_in12[0], w_0545_);
nand (w_0337_, w_0858_, w_0825_);
or (w_0162_, w_0220_, w_0271_);
and (w_0878_, w_0401_, w_0391_);
nand (w_0542_, w_0214_, w_0716_);
xor (w_0518_, new_in18[0], new_in10[0]);
nand (w_0398_, w_0695_, w_0712_);
nand (w_0364_, w_0824_, w_0403_);
nand (w_0444_, w_0858_, w_0495_);
nand (w_0013_, w_0156_, w_0085_);
and (w_0166_, w_0220_, w_0826_);
nand (new_out15[3], w_0396_, w_0151_);
or (w_0944_, w_0564_, w_0290_);
nand (w_0206_, w_0336_, w_0029_);
nand (w_0860_, w_0858_, w_0748_);
nand (w_0759_, w_0695_, w_0499_);
nand (w_0071_, w_0319_, w_0336_);
nand (w_0023_, new_in7[1], w_0824_);
nand (w_0242_, w_0008_, w_0587_);
and (w_0879_, w_0196_, w_0463_);
nand (w_0086_, w_0336_, w_0253_);
nand (w_0082_, w_0022_, w_0618_);
and (w_0322_, w_0409_, w_0775_);
nand (w_0045_, new_in20[0], w_0008_);
xor (w_0746_, w_0706_, w_0509_);
nand (w_0066_, w_0008_, w_0356_);
nand (w_0512_, w_0620_, w_0232_);
nand (w_0304_, new_in8[1], new_in2[1]);
nand (w_0291_, w_0357_, w_0687_);
xor (w_0922_, new_in20[0], w_0452_);
nor (w_0483_, new_in6[0], w_0899_);
nand (w_0870_, w_0254_, w_0642_);
nand (w_0754_, w_0887_, w_0456_);
and (w_0371_, w_0534_, w_0154_);
nand (w_0167_, w_0824_, w_0098_);
nand (w_0792_, w_0008_, w_0732_);
nand (w_0521_, w_0858_, w_0237_);
nand (w_0467_, w_0220_, w_0768_);
xor (w_0835_, w_0202_, w_0784_);
nand (w_0448_, w_0063_, w_0404_);
nand (w_0804_, w_0880_, w_0699_);
and (w_0131_, w_0008_, w_0936_);
xor (w_0367_, new_in19[1], w_0392_);
not (w_0852_, new_in15[1]);
nand (w_0670_, w_0775_, w_0392_);
endmodule
