module new_sub_module1(
    input wire new_in1,
    input wire new_in10,
    input wire new_in11,
    input wire new_in12,
    input wire new_in13,
    input wire new_in14,
    input wire new_in15,
    input wire new_in16,
    input wire new_in2,
    input wire new_in3,
    input wire new_in4,
    input wire new_in5,
    input wire new_in6,
    input wire new_in7,
    input wire new_in8,
    input wire new_in9,
    output wire new_out1,
    output wire new_out10,
    output wire new_out2,
    output wire new_out3,
    output wire new_out4,
    output wire new_out5,
    output wire new_out6,
    output wire new_out7,
    output wire new_out8,
    output wire new_out9
);
wire w_00_;
wire w_01_;
wire w_02_;
wire w_03_;
wire w_04_;
wire w_05_;
wire w_06_;
wire w_07_;
wire w_08_;
wire w_09_;
wire w_10_;
wire w_11_;
wire w_12_;
wire w_13_;
wire w_14_;
wire w_15_;
wire w_16_;
wire w_17_;
wire w_18_;
wire w_19_;
wire w_20_;
wire w_21_;
wire w_22_;
wire w_23_;
wire w_24_;
wire w_25_;
wire w_26_;
wire w_27_;
wire w_28_;
wire w_29_;
wire w_30_;
wire w_31_;
wire w_32_;
wire w_33_;
wire w_34_;
wire w_35_;
wire w_36_;
wire w_37_;
wire w_38_;
wire w_39_;
and (w_37_, new_in9, new_in11);
xor (w_11_, new_in2, w_33_);
xor (w_16_, new_in11, new_in10);
nand (w_14_, new_in7, new_in1);
xor (new_out2, w_10_, w_04_);
and (w_15_, w_31_, w_30_);
and (w_35_, new_in1, new_in16);
xor (new_out7, w_00_, w_36_);
and (new_out1, w_21_, w_01_);
and (w_38_, new_in14, new_in6);
not (w_13_, new_in3);
not (w_21_, w_10_);
nor (w_30_, new_in13, w_23_);
xor (w_28_, w_34_, w_32_);
nor (w_18_, new_in15, w_11_);
nor (w_25_, new_in15, new_in7);
nor (w_23_, new_in6, w_14_);
xor (new_out9, w_18_, w_28_);
xor (w_04_, new_out9, new_out3);
and (w_29_, w_02_, w_25_);
nor (w_39_, w_28_, w_15_);
and (w_33_, new_in4, new_in5);
and (w_06_, w_18_, w_28_);
and (w_34_, w_13_, new_in14);
xor (new_out4, w_18_, w_15_);
and (w_36_, w_06_, w_15_);
and (w_19_, w_22_, w_20_);
not (w_17_, w_03_);
and (w_24_, w_03_, w_39_);
nor (w_32_, new_in12, new_in9);
xor (w_12_, new_in16, new_in8);
xor (w_00_, w_03_, w_10_);
and (w_20_, w_33_, w_38_);
and (w_05_, w_26_, w_29_);
xor (w_10_, w_19_, w_05_);
and (w_01_, w_09_, w_24_);
not (new_out5, w_00_);
xor (new_out10, w_18_, w_00_);
xor (new_out3, w_17_, w_15_);
nor (w_03_, w_16_, w_12_);
nand (w_31_, new_in6, w_14_);
xor (new_out6, w_21_, w_07_);
nor (w_08_, new_in8, new_in10);
xor (w_07_, w_28_, w_15_);
xor (new_out8, w_09_, w_24_);
and (w_26_, w_27_, w_08_);
and (w_22_, w_35_, w_37_);
or (w_09_, new_in15, w_11_);
nor (w_27_, new_in12, new_in2);
nor (w_02_, new_in3, new_in13);
endmodule

module new_sub_module2(
    input wire [5:0] new_in10,
    input wire [5:0] new_in11,
    input wire [5:0] new_in12,
    input wire [5:0] new_in14,
    input wire [5:0] new_in4,
    input wire [5:0] new_in6,
    input wire [5:0] new_in7,
    input wire [5:0] new_in8,
    input wire [7:0] new_in1,
    input wire [7:0] new_in13,
    input wire [7:0] new_in15,
    input wire [7:0] new_in16,
    input wire [7:0] new_in2,
    input wire [7:0] new_in3,
    input wire [7:0] new_in5,
    input wire [7:0] new_in9,
    output wire [5:0] new_out1,
    output wire [5:0] new_out11,
    output wire [5:0] new_out14,
    output wire [5:0] new_out16,
    output wire [5:0] new_out17,
    output wire [5:0] new_out18,
    output wire [5:0] new_out20,
    output wire [5:0] new_out23,
    output wire [5:0] new_out4,
    output wire [5:0] new_out5,
    output wire [5:0] new_out7,
    output wire [5:0] new_out8,
    output wire [7:0] new_out10,
    output wire [7:0] new_out12,
    output wire [7:0] new_out13,
    output wire [7:0] new_out15,
    output wire [7:0] new_out19,
    output wire [7:0] new_out2,
    output wire [7:0] new_out21,
    output wire [7:0] new_out22,
    output wire [7:0] new_out24,
    output wire [7:0] new_out3,
    output wire [7:0] new_out6,
    output wire [7:0] new_out9
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
wire w_0945_;
wire w_0946_;
wire w_0947_;
wire w_0948_;
wire w_0949_;
wire w_0950_;
wire w_0951_;
wire w_0952_;
wire w_0953_;
wire w_0954_;
wire w_0955_;
wire w_0956_;
wire w_0957_;
wire w_0958_;
wire w_0959_;
wire w_0960_;
wire w_0961_;
wire w_0962_;
wire w_0963_;
wire w_0964_;
wire w_0965_;
wire w_0966_;
wire w_0967_;
wire w_0968_;
wire w_0969_;
wire w_0970_;
wire w_0971_;
wire w_0972_;
wire w_0973_;
wire w_0974_;
wire w_0975_;
wire w_0976_;
wire w_0977_;
wire w_0978_;
wire w_0979_;
wire w_0980_;
wire w_0981_;
wire w_0982_;
wire w_0983_;
wire w_0984_;
wire w_0985_;
wire w_0986_;
wire w_0987_;
wire w_0988_;
wire w_0989_;
wire w_0990_;
wire w_0991_;
wire w_0992_;
wire w_0993_;
wire w_0994_;
wire w_0995_;
wire w_0996_;
wire w_0997_;
wire w_0998_;
wire w_0999_;
wire w_1000_;
wire w_1001_;
wire w_1002_;
wire w_1003_;
wire w_1004_;
wire w_1005_;
wire w_1006_;
wire w_1007_;
wire w_1008_;
wire w_1009_;
wire w_1010_;
wire w_1011_;
wire w_1012_;
wire w_1013_;
wire w_1014_;
wire w_1015_;
wire w_1016_;
wire w_1017_;
wire w_1018_;
wire w_1019_;
wire w_1020_;
wire w_1021_;
wire w_1022_;
wire w_1023_;
wire w_1024_;
wire w_1025_;
wire w_1026_;
wire w_1027_;
wire w_1028_;
wire w_1029_;
wire w_1030_;
wire w_1031_;
wire w_1032_;
wire w_1033_;
wire w_1034_;
wire w_1035_;
wire w_1036_;
wire w_1037_;
wire w_1038_;
wire w_1039_;
wire w_1040_;
wire w_1041_;
wire w_1042_;
wire w_1043_;
wire w_1044_;
wire w_1045_;
wire w_1046_;
wire w_1047_;
wire w_1048_;
wire w_1049_;
wire w_1050_;
wire w_1051_;
wire w_1052_;
wire w_1053_;
wire w_1054_;
wire w_1055_;
wire w_1056_;
wire w_1057_;
wire w_1058_;
wire w_1059_;
wire w_1060_;
wire w_1061_;
wire w_1062_;
wire w_1063_;
wire w_1064_;
wire w_1065_;
wire w_1066_;
wire w_1067_;
wire w_1068_;
wire w_1069_;
wire w_1070_;
wire w_1071_;
wire w_1072_;
wire w_1073_;
wire w_1074_;
wire w_1075_;
wire w_1076_;
wire w_1077_;
wire w_1078_;
wire w_1079_;
wire w_1080_;
wire w_1081_;
wire w_1082_;
wire w_1083_;
wire w_1084_;
wire w_1085_;
wire w_1086_;
wire w_1087_;
wire w_1088_;
wire w_1089_;
wire w_1090_;
wire w_1091_;
wire w_1092_;
wire w_1093_;
wire w_1094_;
wire w_1095_;
wire w_1096_;
wire w_1097_;
wire w_1098_;
wire w_1099_;
wire w_1100_;
wire w_1101_;
wire w_1102_;
wire w_1103_;
wire w_1104_;
wire w_1105_;
wire w_1106_;
wire w_1107_;
wire w_1108_;
wire w_1109_;
wire w_1110_;
wire w_1111_;
wire w_1112_;
wire w_1113_;
wire w_1114_;
wire w_1115_;
wire w_1116_;
wire w_1117_;
wire w_1118_;
wire w_1119_;
wire w_1120_;
wire w_1121_;
wire w_1122_;
wire w_1123_;
wire w_1124_;
wire w_1125_;
wire w_1126_;
wire w_1127_;
wire w_1128_;
wire w_1129_;
wire w_1130_;
wire w_1131_;
wire w_1132_;
wire w_1133_;
wire w_1134_;
wire w_1135_;
wire w_1136_;
wire w_1137_;
wire w_1138_;
wire w_1139_;
wire w_1140_;
wire w_1141_;
wire w_1142_;
wire w_1143_;
wire w_1144_;
wire w_1145_;
wire w_1146_;
wire w_1147_;
wire w_1148_;
wire w_1149_;
wire w_1150_;
wire w_1151_;
wire w_1152_;
wire w_1153_;
wire w_1154_;
wire w_1155_;
wire w_1156_;
wire w_1157_;
wire w_1158_;
wire w_1159_;
wire w_1160_;
wire w_1161_;
wire w_1162_;
wire w_1163_;
wire w_1164_;
wire w_1165_;
wire w_1166_;
wire w_1167_;
wire w_1168_;
wire w_1169_;
wire w_1170_;
wire w_1171_;
wire w_1172_;
wire w_1173_;
wire w_1174_;
wire w_1175_;
wire w_1176_;
wire w_1177_;
wire w_1178_;
wire w_1179_;
wire w_1180_;
wire w_1181_;
wire w_1182_;
wire w_1183_;
wire w_1184_;
wire w_1185_;
wire w_1186_;
wire w_1187_;
wire w_1188_;
wire w_1189_;
wire w_1190_;
wire w_1191_;
wire w_1192_;
wire w_1193_;
wire w_1194_;
wire w_1195_;
wire w_1196_;
wire w_1197_;
wire w_1198_;
wire w_1199_;
wire w_1200_;
wire w_1201_;
wire w_1202_;
wire w_1203_;
wire w_1204_;
wire w_1205_;
wire w_1206_;
wire w_1207_;
wire w_1208_;
wire w_1209_;
wire w_1210_;
wire w_1211_;
wire w_1212_;
wire w_1213_;
wire w_1214_;
wire w_1215_;
wire w_1216_;
wire w_1217_;
wire w_1218_;
wire w_1219_;
wire w_1220_;
wire w_1221_;
wire w_1222_;
wire w_1223_;
wire w_1224_;
wire w_1225_;
wire w_1226_;
wire w_1227_;
wire w_1228_;
wire w_1229_;
wire w_1230_;
xor (w_1199_, w_0765_, w_0777_);
xor (w_0349_, w_0444_, w_0341_);
xor (w_0147_, w_1140_, w_0366_);
xor (w_0669_, w_0052_, w_0698_);
nand (w_0157_, w_0780_, w_0827_);
nand (w_0877_, w_1064_, w_0241_);
xor (new_out1[4], w_0057_, w_1030_);
nand (w_0396_, new_in13[4], w_0778_);
and (w_0923_, w_1009_, w_0248_);
and (w_1070_, w_0490_, w_0479_);
nand (w_1001_, w_0810_, w_0373_);
nand (w_0567_, w_0415_, w_1119_);
or (new_out15[7], w_0857_, w_1141_);
and (w_0208_, w_0153_, w_0145_);
xor (w_0588_, w_0967_, w_0751_);
or (w_0388_, w_0841_, w_0422_);
nand (w_0135_, w_0199_, w_1007_);
xor (w_0428_, new_in13[6], w_0344_);
nand (w_0693_, new_in16[3], new_in3[3]);
xor (w_1119_, w_0500_, w_1049_);
xor (w_0212_, w_0351_, w_0969_);
xor (w_0219_, w_1001_, w_0727_);
xor (w_0870_, w_0999_, w_0386_);
xor (new_out11[3], w_0776_, w_0835_);
nand (w_0487_, w_0606_, w_1220_);
or (new_out15[1], w_0436_, w_0785_);
xor (w_0880_, new_in6[0], w_1206_);
nand (w_1158_, w_0620_, w_1095_);
nand (w_0667_, w_0356_, w_0238_);
and (w_0760_, new_in3[0], new_in16[0]);
and (w_0781_, w_0097_, w_0878_);
xor (w_0843_, new_in14[0], new_in6[1]);
or (w_0559_, w_0394_, w_1112_);
and (w_0689_, new_in5[0], w_0756_);
or (w_0960_, w_0642_, w_0463_);
nand (w_0823_, w_0170_, w_0439_);
nand (w_0527_, w_0087_, w_0435_);
nand (w_0924_, w_0207_, w_0753_);
nand (w_0330_, new_in16[4], new_in3[4]);
xor (w_1066_, w_1052_, w_0501_);
nand (w_0498_, w_0451_, w_1216_);
nand (w_0400_, w_1097_, w_0027_);
xor (w_0307_, w_0076_, w_0939_);
xor (w_0698_, new_in11[1], w_0271_);
or (w_0680_, w_0675_, w_1171_);
xor (w_0532_, w_0606_, w_0155_);
nand (w_0086_, w_0596_, w_0376_);
xor (w_0055_, w_0193_, w_0978_);
nand (w_0953_, w_0235_, w_0918_);
and (w_0181_, w_0590_, w_0091_);
xor (w_0623_, w_1224_, w_1147_);
nand (w_0080_, w_0545_, new_out8[4]);
nand (w_0293_, new_in11[1], w_0271_);
xor (new_out11[1], w_0119_, w_0382_);
xor (new_out23[2], w_1048_, w_0686_);
or (w_0742_, w_0298_, w_1015_);
xor (w_0981_, new_in6[5], w_0115_);
xor (w_0701_, w_1197_, w_0551_);
nand (w_0574_, new_in14[4], w_0865_);
nand (w_0297_, w_0433_, w_1041_);
or (w_0685_, w_0449_, w_0107_);
nand (w_0415_, w_0998_, w_0014_);
xor (w_0426_, w_1155_, w_0980_);
nand (w_0971_, w_1155_, w_0980_);
nand (w_1215_, w_0531_, w_1129_);
and (w_0751_, w_0621_, w_1108_);
nand (w_0286_, new_in1[5], w_0480_);
xor (w_1153_, new_in13[1], w_0156_);
xor (w_0514_, w_1137_, w_0456_);
xor (w_0048_, new_in11[0], w_0651_);
nand (w_0238_, w_0314_, w_0218_);
not (new_out19[6], w_0027_);
nand (w_1081_, new_in10[5], w_0413_);
or (w_0738_, w_0707_, w_0367_);
xor (w_0422_, w_0856_, w_0903_);
and (w_0235_, w_0006_, w_0414_);
nor (w_0868_, w_0444_, w_0341_);
xor (w_0156_, w_0536_, w_0550_);
xor (new_out7[0], w_0205_, w_0246_);
nand (w_0754_, w_0039_, w_0340_);
xor (new_out12[2], w_1037_, w_0448_);
not (w_0743_, w_0107_);
xor (new_out21[7], w_0284_, w_1021_);
and (new_out13[0], w_0670_, w_0738_);
nand (w_1089_, w_0930_, w_0094_);
xor (new_out12[5], w_1220_, w_1012_);
xor (w_0713_, new_in5[4], w_0704_);
xor (w_0907_, w_1113_, w_0395_);
xor (w_1213_, new_in14[5], w_0645_);
xor (w_0439_, w_0785_, w_0673_);
nand (w_0979_, w_1187_, w_0080_);
xor (w_0969_, w_1155_, w_0038_);
nand (w_0986_, w_0718_, w_0478_);
xor (w_0459_, w_1140_, w_0021_);
xor (new_out7[1], w_1212_, w_0138_);
xor (w_0581_, new_in9[5], new_in13[5]);
xor (w_0007_, w_0866_, w_0914_);
and (w_0028_, w_1140_, w_0490_);
nand (w_0832_, new_in12[1], w_0148_);
nand (w_0836_, w_0791_, w_1145_);
nand (w_0842_, w_0699_, w_1038_);
xor (w_0231_, w_0038_, w_0020_);
nand (w_0195_, w_0992_, w_0981_);
not (w_0639_, w_0720_);
xor (w_0927_, w_1071_, w_0349_);
xor (w_1048_, w_1128_, w_1205_);
nand (w_0859_, new_in2[1], w_0405_);
nand (new_out3[4], w_0592_, w_0904_);
xor (w_0001_, w_0267_, w_0244_);
nand (w_0253_, w_0332_, w_1126_);
xor (new_out21[6], w_0098_, w_0732_);
nand (w_0243_, w_0017_, w_0383_);
xor (w_0013_, w_1105_, w_0663_);
nand (w_1118_, w_1003_, w_0936_);
xor (new_out20[1], w_1097_, w_0027_);
nand (w_1023_, new_in6[1], w_1014_);
not (w_0758_, w_1133_);
nand (w_0892_, w_0506_, w_1047_);
xor (w_0044_, new_in14[2], w_0768_);
nand (w_0408_, w_0038_, w_1071_);
nand (w_0417_, w_0589_, w_0133_);
nor (w_0202_, w_1140_, w_0707_);
xor (w_0939_, new_in12[2], w_0870_);
nand (w_0485_, w_0016_, w_0171_);
nand (w_0136_, new_in8[2], new_in7[2]);
or (w_0956_, new_in13[3], w_0850_);
nand (w_1052_, w_0390_, w_1051_);
xor (w_0974_, w_0076_, w_0120_);
xor (w_0436_, w_0948_, w_0763_);
xor (w_0138_, w_0673_, w_1205_);
nand (w_0564_, w_1110_, w_0944_);
nand (w_0573_, w_0638_, w_0660_);
xor (w_0662_, w_0126_, w_0418_);
xor (w_0525_, w_0228_, w_1071_);
xor (w_0651_, new_in8[1], new_in7[0]);
xor (w_0036_, w_0122_, w_0571_);
nand (w_1187_, w_0907_, w_1133_);
xor (w_0370_, new_in1[0], w_0427_);
xor (w_0825_, w_0182_, w_0438_);
xor (w_0217_, new_in15[4], w_0687_);
nand (w_0886_, w_0654_, w_0706_);
nand (w_0716_, w_0431_, w_0721_);
xor (w_0943_, w_1226_, w_0855_);
xor (w_0403_, w_1227_, w_0796_);
xor (w_0082_, new_in11[2], w_0036_);
xor (w_0483_, w_0074_, w_0246_);
xor (w_0079_, w_0599_, w_0049_);
nand (w_0622_, w_1121_, w_0877_);
nand (w_0247_, w_0924_, w_0745_);
xor (new_out18[5], w_0305_, w_0837_);
nand (w_0336_, w_0125_, w_0441_);
xor (new_out10[4], w_0298_, w_1015_);
xor (w_1190_, w_0678_, w_0966_);
nand (w_0008_, w_0530_, w_0703_);
xor (w_0753_, w_0415_, w_1119_);
xor (w_1105_, w_0845_, w_0840_);
xor (w_0613_, w_0634_, w_0580_);
nand (w_0469_, w_0482_, w_1122_);
nand (w_0442_, w_1166_, w_0393_);
nand (w_0420_, w_0437_, w_0306_);
xor (w_0094_, new_in1[5], new_in15[5]);
xor (w_1080_, w_0343_, w_0428_);
and (w_0256_, w_1137_, w_0456_);
xor (new_out22[7], w_0952_, w_0123_);
nand (w_0472_, w_0152_, w_0678_);
nand (w_1221_, w_0941_, w_0389_);
nand (w_0518_, new_in9[5], new_in13[5]);
and (w_0394_, w_1019_, w_1157_);
nand (w_0784_, new_in5[6], w_0011_);
nand (w_0014_, w_0692_, w_1165_);
xor (w_1164_, new_in15[5], w_0748_);
xor (w_1138_, w_0474_, w_0277_);
and (w_1033_, w_0589_, w_0522_);
xor (w_0722_, w_0102_, w_0255_);
xor (w_0770_, new_out2[0], w_0367_);
xor (w_1014_, w_0994_, w_0867_);
and (w_0611_, w_0408_, w_0275_);
nand (w_0348_, w_0267_, w_0244_);
nand (w_0132_, new_in8[5], new_in7[5]);
nand (w_0750_, w_1010_, w_1071_);
not (w_1043_, new_in4[0]);
nand (w_0249_, w_0760_, w_1115_);
nand (w_0056_, new_in5[2], w_0128_);
xor (w_0947_, w_0620_, w_0367_);
xor (w_0445_, w_0718_, w_0478_);
or (w_0441_, w_1105_, w_0615_);
xor (w_0179_, w_0180_, w_1195_);
nand (w_0104_, w_0452_, w_0310_);
xor (w_0530_, w_1010_, w_1071_);
xor (new_out21[5], w_0345_, w_1099_);
xor (w_0023_, new_in2[4], w_0509_);
xor (w_0174_, w_0908_, w_1033_);
nand (w_0017_, w_0213_, w_0081_);
nand (w_0373_, w_0002_, w_1016_);
nand (w_0978_, w_0118_, w_0680_);
or (w_1108_, new_in9[6], new_in13[6]);
xor (w_0752_, w_1037_, w_1133_);
xor (w_1205_, w_1037_, w_1105_);
xor (new_out5[5], w_0666_, w_0224_);
nand (w_0236_, w_0040_, w_0328_);
nand (w_0796_, w_0396_, w_0100_);
nand (w_0275_, w_0494_, w_1184_);
nand (w_0961_, w_1168_, w_1004_);
xor (w_1037_, w_0654_, w_0706_);
xor (w_0802_, new_in2[7], w_0457_);
or (w_0890_, w_0758_, w_0449_);
nand (w_0546_, new_in12[3], w_0849_);
xor (new_out20[5], w_0829_, w_0813_);
nand (w_1168_, new_in10[4], w_0001_);
nand (w_0437_, new_in1[2], w_0007_);
nand (w_0854_, w_0635_, w_1044_);
xor (w_0650_, new_in3[0], new_in16[0]);
and (w_0423_, w_0750_, w_0130_);
and (w_0298_, w_0312_, w_0033_);
xor (w_0671_, w_1210_, w_0226_);
not (w_1203_, w_0024_);
and (w_1195_, w_0841_, w_0856_);
xor (w_0786_, w_1009_, w_0079_);
xor (w_0645_, w_0961_, w_0729_);
xor (w_0414_, w_0902_, w_0864_);
not (w_0260_, w_0678_);
xor (w_0856_, new_in9[0], w_0830_);
nand (w_0343_, w_0464_, w_1067_);
xor (new_out10[0], w_1140_, w_0490_);
xor (w_0061_, new_in8[3], new_in7[2]);
xor (new_out5[3], w_0858_, new_out13[5]);
nand (w_0184_, w_1158_, w_0124_);
and (w_0331_, w_1069_, w_0622_);
nand (w_0322_, w_0258_, new_out8[2]);
nand (w_0434_, w_0419_, w_1156_);
not (w_0380_, new_out2[0]);
xor (new_out8[1], w_0436_, w_0673_);
nand (w_0201_, w_0351_, w_0969_);
and (w_0198_, new_out8[0], w_1140_);
xor (new_out22[1], w_1151_, w_0352_);
xor (w_0777_, w_1124_, w_0836_);
nand (w_0190_, w_0157_, w_0053_);
nand (w_0000_, w_1093_, w_0893_);
and (w_0092_, new_in6[0], w_1206_);
xor (w_0871_, w_0339_, w_0786_);
xor (w_0034_, w_0494_, w_1184_);
nand (w_0885_, w_1228_, w_0261_);
nand (w_0458_, w_0738_, w_0828_);
and (w_0812_, w_0412_, w_0046_);
nand (w_0497_, new_in1[1], w_1056_);
xor (w_0830_, new_in13[0], w_0370_);
and (new_out6[3], w_0020_, w_0927_);
xor (w_0542_, w_1220_, w_0806_);
nand (w_0711_, w_1162_, w_0288_);
not (w_1135_, w_0398_);
xor (w_1022_, w_0711_, w_0883_);
nand (w_1196_, new_in3[2], new_in16[2]);
nand (w_1078_, w_0151_, w_1091_);
nand (w_0419_, w_0178_, w_0313_);
xor (w_0595_, w_0449_, w_0743_);
xor (w_1123_, w_0325_, w_0853_);
nand (w_1028_, new_in5[5], w_0189_);
xor (new_out24[0], w_0380_, new_out10[0]);
nand (w_0215_, w_0047_, w_0581_);
xor (new_out21[1], w_0709_, w_0443_);
xor (new_out14[4], w_0678_, w_0106_);
and (w_1059_, w_1176_, w_0533_);
xor (w_0261_, new_in15[7], w_0943_);
xor (w_1084_, w_0017_, w_0383_);
xor (w_0997_, w_0363_, w_0499_);
xor (new_out10[2], w_1024_, w_0724_);
or (w_0762_, w_1225_, w_1059_);
nand (new_out3[6], w_0246_, w_0746_);
nand (w_1110_, w_0694_, w_0314_);
xor (w_0789_, w_0696_, w_0422_);
nand (w_1051_, w_0102_, w_0255_);
and (w_0371_, new_in9[3], new_in13[3]);
or (w_0506_, w_1147_, w_0245_);
xor (w_1200_, w_1085_, w_1159_);
xor (w_0031_, w_0655_, w_0231_);
nand (w_0826_, w_1076_, w_0239_);
xor (new_out5[4], w_0303_, w_0168_);
nand (w_0097_, w_1178_, w_0259_);
and (w_0332_, w_0276_, w_0749_);
nand (w_0808_, new_in15[2], w_0899_);
not (w_0879_, w_0141_);
xor (w_0864_, w_0638_, w_0660_);
xor (w_0143_, w_0307_, w_0230_);
xor (w_0096_, new_in1[3], w_1132_);
nand (w_0691_, w_0090_, w_0947_);
xor (new_out22[5], w_0934_, w_0263_);
nand (w_1004_, w_1079_, w_0468_);
xor (w_0576_, w_0431_, w_0721_);
xor (w_0435_, new_in12[3], w_0849_);
nand (w_0199_, new_in15[4], w_0687_);
nand (w_0894_, w_0994_, w_0867_);
xor (w_1194_, new_in10[0], w_0769_);
nand (w_0375_, w_1073_, w_0225_);
xor (w_0281_, new_in6[5], new_in14[4]);
xor (w_1147_, w_1008_, w_0719_);
nand (w_0193_, w_0132_, w_0643_);
xor (w_0606_, w_0172_, w_0681_);
xor (w_0491_, w_0399_, w_0655_);
nand (w_0995_, w_1229_, w_0315_);
xor (w_0676_, w_1221_, w_0217_);
xor (w_0747_, w_0060_, w_0641_);
and (w_0990_, w_0153_, w_1214_);
xor (w_0898_, new_in9[4], new_in13[4]);
xor (w_0405_, w_0760_, w_1115_);
xor (w_0493_, w_0625_, w_0891_);
nand (w_0658_, w_0076_, w_1037_);
nand (w_1029_, w_0182_, w_0438_);
xor (w_1149_, w_0172_, w_0305_);
xor (w_0790_, w_0397_, w_0604_);
and (w_0406_, w_1220_, w_0806_);
xor (w_0901_, w_0258_, new_out8[2]);
and (w_0489_, w_1177_, w_0400_);
nand (w_0929_, w_0608_, w_0804_);
nand (w_1091_, w_0942_, w_0539_);
nand (w_0977_, w_0523_, w_0957_);
nand (w_0192_, new_in9[4], new_in13[4]);
xor (w_0571_, new_in8[2], new_in7[2]);
xor (w_0795_, w_0152_, w_0678_);
nand (w_0374_, w_0505_, w_0755_);
xor (w_1143_, w_0649_, w_0636_);
nand (w_0715_, w_0961_, w_0729_);
and (w_0934_, w_0150_, w_0985_);
nand (w_0196_, w_1013_, w_1199_);
xor (w_0834_, new_in1[2], w_0007_);
nand (w_0062_, w_0030_, w_1018_);
nand (w_1219_, w_0832_, w_0166_);
xor (w_0386_, new_in6[2], new_in14[1]);
nand (w_0121_, w_0984_, w_0973_);
or (w_0819_, w_0991_, w_1183_);
nand (w_0670_, w_0707_, w_0367_);
nand (w_0258_, w_0142_, w_0736_);
nand (w_0496_, w_0020_, w_0837_);
nand (w_0225_, w_0987_, w_0431_);
xor (w_0185_, new_in8[4], new_in7[4]);
nand (w_1216_, w_0168_, w_1082_);
nand (w_0726_, w_0623_, w_0034_);
xor (w_0778_, w_0485_, w_0242_);
nand (w_1061_, w_1009_, w_0079_);
and (new_out17[5], w_0623_, w_1128_);
xor (new_out14[0], w_0074_, w_0147_);
xor (w_0120_, w_1219_, w_0495_);
xor (w_0916_, w_0021_, w_0500_);
nand (new_out3[7], w_0041_, w_1205_);
nand (w_0549_, w_0119_, w_0382_);
nand (w_0630_, w_0222_, w_1074_);
nand (w_0019_, w_0175_, w_1110_);
xor (w_0558_, w_0431_, w_0467_);
xor (w_1092_, new_in5[0], w_0756_);
nand (w_0087_, w_0647_, w_1020_);
xor (w_0592_, w_0857_, w_0152_);
xor (w_0959_, w_1011_, w_0004_);
not (w_1090_, new_in2[7]);
nand (w_0872_, w_0859_, w_0018_);
and (w_1136_, w_0404_, w_0210_);
xor (new_out13[4], w_1161_, w_0875_);
and (w_0220_, w_0824_, w_0644_);
xor (w_0490_, w_0718_, w_0759_);
xor (w_0020_, w_0087_, w_0435_);
nand (w_1058_, w_0967_, w_1108_);
nand (w_0102_, w_0358_, w_1131_);
nand (w_0565_, w_0250_, w_0445_);
xor (w_0840_, new_in5[1], w_0273_);
nand (w_0920_, new_in13[3], w_0850_);
nand (w_0058_, w_1118_, w_1140_);
xor (new_out12[7], w_0926_, w_1185_);
or (w_0444_, w_1017_, w_0674_);
not (w_0425_, w_0606_);
nand (w_1142_, w_0083_, w_0544_);
nand (w_1064_, w_1037_, w_0848_);
nand (w_0503_, w_1023_, w_0653_);
nand (w_1063_, w_0237_, w_0015_);
nand (w_0824_, w_0229_, w_0134_);
nand (w_0402_, w_0603_, w_0305_);
xor (w_1159_, new_in12[4], w_0219_);
nand (w_0695_, new_in2[7], w_1066_);
xor (w_1181_, new_in16[4], new_in3[4]);
nand (w_0356_, w_0203_, w_0819_);
xor (w_0857_, w_1225_, w_1059_);
xor (w_0794_, w_0689_, w_0628_);
nand (w_0608_, w_0678_, w_0966_);
nand (w_1217_, w_0502_, w_0063_);
nand (w_0683_, w_0621_, w_1058_);
nand (w_0589_, new_in8[3], new_in7[3]);
nand (w_1192_, new_in1[4], w_0676_);
and (w_0876_, w_0726_, w_0022_);
xor (w_0629_, w_0927_, w_0075_);
nand (w_0998_, w_0592_, w_1230_);
xor (new_out10[5], new_out23[0], w_0429_);
and (w_0067_, w_0547_, w_0757_);
nand (w_0593_, w_1212_, w_0138_);
xor (w_0323_, w_0074_, w_0211_);
nand (w_0279_, w_0652_, w_0922_);
xor (new_out10[6], w_0232_, w_0483_);
nand (w_1125_, w_0730_, w_0932_);
nand (w_1204_, w_0013_, w_0958_);
nand (w_0757_, w_0765_, w_0777_);
nand (w_0725_, w_0246_, w_0424_);
nand (w_0040_, w_0402_, w_0773_);
xor (w_0853_, w_0502_, w_0063_);
nand (w_0390_, new_in16[6], new_in3[6]);
not (w_0085_, w_0642_);
not (w_1010_, w_0038_);
nand (w_1179_, w_0240_, w_0713_);
xor (w_0134_, w_0168_, w_0059_);
nand (w_0440_, w_0385_, w_0086_);
or (w_1156_, w_0181_, w_0906_);
and (w_1151_, w_0707_, w_0770_);
nand (w_0547_, w_1124_, w_0836_);
nand (w_0167_, w_0689_, w_0628_);
xor (w_0463_, new_in1[3], new_in15[3]);
xor (w_1175_, new_in4[5], w_0800_);
nand (w_1155_, w_0733_, w_0421_);
nand (w_0922_, w_1024_, w_0724_);
xor (w_1230_, w_0545_, new_out8[4]);
nand (w_1011_, w_0983_, w_0320_);
xor (w_1049_, new_out8[5], w_0979_);
xor (new_out12[3], w_0694_, w_1209_);
nand (w_1041_, w_0473_, w_0691_);
xor (w_0642_, w_0484_, w_0308_);
xor (w_1227_, new_in13[5], w_1057_);
nand (w_0233_, w_0074_, w_0246_);
nand (w_0933_, new_in2[3], w_0790_);
nand (w_0599_, w_1089_, w_0762_);
xor (w_1032_, new_in2[4], w_0556_);
nand (w_1139_, w_0025_, w_0553_);
xor (w_1057_, w_0635_, w_1044_);
xor (w_1034_, new_in9[3], w_0671_);
not (w_0666_, new_out13[7]);
xor (new_out14[2], w_0707_, w_0488_);
nand (w_0539_, w_1106_, w_0782_);
xor (w_0641_, w_0404_, w_0210_);
nand (w_0145_, w_0587_, w_1214_);
nand (w_0316_, w_0842_, w_0471_);
nand (new_out3[3], w_0655_, w_0459_);
xor (new_out21[2], w_0664_, w_1053_);
or (w_0232_, w_0833_, w_0309_);
xor (new_out13[2], w_0260_, w_0449_);
xor (w_0900_, new_in14[4], w_0865_);
nand (w_1208_, new_in1[7], w_1170_);
xor (w_0159_, w_0995_, w_0646_);
xor (w_0257_, w_0580_, w_0901_);
nand (w_0553_, w_0398_, w_0789_);
xor (w_0467_, w_0276_, w_0749_);
xor (w_0649_, new_in5[3], w_1222_);
xor (w_0855_, new_in5[7], w_0364_);
nand (w_0030_, w_1086_, w_0657_);
xor (w_0740_, w_1224_, w_0681_);
xor (new_out12[1], w_0038_, w_0475_);
nand (w_0346_, w_0634_, w_0580_);
or (w_1109_, w_0554_, w_0551_);
nand (w_0618_, w_1040_, w_0740_);
not (w_0999_, new_in4[1]);
xor (w_0838_, w_0207_, w_0753_);
and (w_0874_, w_0971_, w_0543_);
nand (w_0967_, w_0518_, w_0215_);
xor (new_out2[5], w_0895_, w_0892_);
nand (w_0053_, w_1070_, w_0563_);
xor (new_out11[2], w_0640_, w_0613_);
not (w_0993_, w_0139_);
xor (w_0600_, w_0500_, w_0158_);
nand (w_0351_, w_1061_, w_0862_);
nand (w_0946_, new_in4[4], w_0317_);
xor (w_0254_, new_in5[2], w_0128_);
nand (w_0745_, w_0838_, w_0434_);
nand (w_0391_, w_1215_, w_0601_);
xor (new_out13[7], w_0606_, w_1141_);
xor (new_out14[5], w_0837_, w_0600_);
nand (w_0569_, new_in8[1], new_in7[1]);
nand (w_1002_, w_0450_, w_0411_);
xor (w_0597_, new_in2[1], w_0405_);
nand (w_1188_, w_0000_, w_0441_);
and (w_0991_, w_0065_, w_0200_);
xor (w_0341_, new_in12[5], w_0861_);
xor (w_0172_, w_0121_, w_0928_);
nand (w_0237_, w_0697_, w_0108_);
xor (w_1056_, w_0117_, w_1027_);
not (w_0603_, w_0172_);
and (w_0119_, w_1140_, w_0431_);
or (w_0962_, w_0325_, w_0853_);
xor (w_0168_, w_0598_, w_0456_);
xor (w_0460_, w_0596_, w_0376_);
xor (w_0509_, new_in3[0], new_in16[4]);
and (w_0161_, w_0515_, w_0960_);
xor (w_0702_, w_0598_, w_0406_);
xor (w_0987_, w_0169_, w_0988_);
xor (new_out2[6], w_0168_, w_1082_);
xor (new_out22[3], w_1036_, w_0929_);
and (w_1144_, new_in13[0], w_0370_);
xor (w_0411_, w_0246_, w_0424_);
nand (w_0626_, w_1140_, w_0020_);
nand (w_0486_, w_0349_, w_0456_);
nor (w_1099_, w_0500_, w_0615_);
not (w_0528_, w_1161_);
or (new_out15[4], w_0907_, w_0528_);
nand (w_0958_, w_0568_, w_1152_);
nand (w_0311_, w_0125_, w_1188_);
nand (w_0881_, w_0970_, w_0249_);
xor (new_out21[4], w_0278_, w_0338_);
nand (w_0621_, new_in9[6], new_in13[6]);
xor (w_0430_, w_0907_, w_1198_);
nand (w_1006_, w_0051_, w_0820_);
xor (w_0895_, w_0606_, w_1220_);
xor (w_0418_, new_in14[2], new_in6[3]);
nand (w_0327_, w_0866_, w_0914_);
not (w_0775_, w_0857_);
xor (new_out24[2], w_0107_, new_out10[2]);
not (w_0245_, w_0229_);
xor (new_out7[4], w_0208_, w_0583_);
nand (w_0453_, w_0329_, w_0362_);
xor (w_0148_, w_0083_, w_0544_);
nand (w_0473_, w_0620_, w_0367_);
nand (w_0610_, new_in11[3], w_0174_);
not (w_0945_, w_0034_);
nand (w_0952_, w_0851_, w_1050_);
xor (w_0548_, w_1135_, w_0789_);
nand (w_0637_, w_0552_, w_0667_);
nand (w_0078_, w_0233_, w_1045_);
xor (w_0479_, new_out8[0], w_1140_);
nand (w_0535_, w_0197_, w_1123_);
xor (w_0705_, w_0342_, w_0597_);
or (w_0015_, w_1113_, w_0395_);
and (w_0675_, w_0937_, w_0348_);
nand (w_0792_, w_0416_, w_0099_);
and (w_1148_, w_0735_, w_0921_);
nand (w_0736_, w_0672_, new_out8[1]);
xor (w_0884_, w_0387_, w_0570_);
nand (w_0006_, w_0378_, w_0885_);
xor (w_0382_, w_0907_, w_1224_);
nand (w_0499_, w_1068_, w_0201_);
or (new_out15[3], w_1140_, w_0837_);
xor (w_0555_, w_1144_, w_1153_);
nand (w_0069_, w_0085_, w_0907_);
nand (w_0129_, new_out13[1], w_0803_);
or (w_1146_, w_1071_, w_0655_);
or (w_1094_, new_out10[4], w_0304_);
xor (w_0821_, w_0143_, w_0807_);
xor (w_0302_, w_0047_, w_0581_);
xor (w_1207_, new_in10[4], w_0470_);
or (w_0065_, w_0665_, w_0075_);
nand (w_0776_, w_0346_, w_0465_);
xor (w_0223_, new_in4[0], w_0880_);
and (w_1184_, w_0079_, w_0634_);
nand (w_0016_, new_in1[3], w_1132_);
nand (w_0511_, new_in11[2], w_0036_);
nand (w_1145_, w_1046_, w_0055_);
xor (w_0255_, new_in16[6], new_in3[6]);
xor (w_0326_, w_0447_, w_0296_);
not (w_0295_, w_1155_);
nand (w_0451_, w_0598_, w_0456_);
xor (new_out23[3], new_out13[0], w_0828_);
xor (w_0248_, new_in12[0], w_0223_);
xor (new_out8[4], w_0907_, w_1133_);
nand (w_1054_, new_in10[3], w_0688_);
xor (w_0914_, new_in15[2], w_0899_);
xor (new_out7[2], w_1180_, w_0616_);
nand (w_0194_, w_0890_, w_0071_);
nand (w_0970_, new_in3[1], new_in16[1]);
nand (w_0568_, w_1133_, w_1200_);
or (w_0773_, w_1149_, w_0737_);
xor (new_out23[4], new_out13[1], w_0803_);
xor (w_0234_, w_0356_, w_0109_);
xor (w_0271_, w_0051_, w_0820_);
nand (w_0066_, w_0615_, w_0289_);
nand (w_1223_, w_0895_, w_0892_);
xor (w_0471_, new_in10[3], w_0688_);
or (w_0602_, w_1155_, w_0251_);
nand (w_0358_, new_in16[5], new_in3[5]);
xor (w_0861_, w_0712_, w_0281_);
nand (w_0932_, w_0511_, w_0624_);
nand (w_0088_, w_0057_, w_1030_);
nand (w_1005_, new_out8[5], w_0979_);
or (w_0227_, w_0188_, w_0886_);
or (w_1186_, w_0041_, w_0915_);
nand (w_0300_, w_0497_, w_1026_);
xor (w_0379_, new_in1[6], w_1022_);
xor (new_out8[3], w_1140_, w_0020_);
xor (w_0845_, new_in10[2], w_0101_);
xor (w_0746_, w_0987_, w_0456_);
nand (w_0659_, new_in4[1], w_0873_);
xor (w_0570_, w_1048_, w_0003_);
nand (w_0799_, w_0440_, w_0900_);
nand (w_0940_, w_0066_, w_1150_);
xor (w_1062_, w_0982_, w_1175_);
xor (w_0413_, w_0675_, w_1171_);
xor (w_0163_, w_0079_, w_0152_);
nand (w_1193_, new_in14[1], w_0714_);
nand (w_0783_, new_in6[4], w_0632_);
xor (w_0687_, w_0240_, w_0713_);
xor (w_0566_, w_1161_, w_0561_);
xor (w_0164_, w_1133_, w_1161_);
nand (w_0291_, new_in6[5], w_0115_);
not (w_0625_, new_in4[3]);
not (w_1173_, w_1040_);
nand (w_0222_, new_in12[4], w_0219_);
xor (new_out13[5], w_0021_, w_0615_);
nand (w_0404_, w_1208_, w_0977_);
nand (w_0533_, w_0169_, w_0988_);
nand (w_1067_, w_1227_, w_0796_);
and (w_0042_, new_in10[0], w_0769_);
nand (w_0798_, w_0780_, w_1205_);
xor (w_0364_, w_0394_, w_1112_);
xor (w_0909_, w_1043_, w_0843_);
nand (w_0481_, w_0744_, w_0010_);
xor (new_out1[2], w_0090_, w_0947_);
nand (w_1189_, w_1039_, w_0105_);
and (w_0361_, w_0948_, w_0763_);
xor (w_0561_, w_0991_, w_1183_);
xor (w_1112_, w_1090_, w_1066_);
nand (w_0660_, w_0695_, w_0559_);
nand (w_0504_, w_1042_, w_1181_);
nand (w_0290_, w_1193_, w_0894_);
xor (w_1012_, w_0000_, w_0336_);
xor (new_out5[1], new_out13[3], w_0019_);
nand (w_1229_, new_in13[1], w_0156_);
nand (w_0024_, w_0888_, w_1204_);
xor (w_0492_, w_0041_, w_0915_);
xor (w_0012_, new_in5[0], w_0023_);
xor (w_0111_, w_0923_, w_1155_);
nand (w_0252_, new_in9[1], w_0555_);
not (w_0178_, w_0186_);
nand (w_0464_, new_in13[5], w_1057_);
xor (w_0896_, new_in15[4], new_in1[4]);
xor (w_1134_, w_0305_, w_0606_);
nand (w_0455_, w_0024_, w_0558_);
nand (w_0450_, w_0731_, w_0567_);
xor (w_1035_, new_in7[4], new_in8[5]);
or (w_0905_, w_0180_, w_1195_);
xor (w_0480_, w_1164_, w_0135_);
xor (w_0377_, w_0449_, w_0829_);
nand (w_1160_, w_0996_, w_1117_);
and (new_out17[0], w_0592_, w_0620_);
xor (w_0519_, w_0229_, w_0134_);
or (w_0985_, w_1167_, w_0566_);
xor (w_0158_, w_0143_, w_0964_);
xor (new_out2[7], w_0224_, w_0498_);
xor (w_0478_, new_in1[7], new_in15[7]);
nand (w_0022_, w_1120_, w_1172_);
xor (w_0848_, w_0853_, w_1200_);
xor (w_0495_, new_in12[2], w_0384_);
xor (w_0891_, new_in6[4], new_in14[3]);
nand (w_1074_, w_1085_, w_1159_);
xor (w_0601_, new_in13[7], w_0154_);
xor (w_0011_, w_1078_, w_0524_);
nand (w_0100_, w_0474_, w_0277_);
xor (w_0149_, new_in11[2], w_0061_);
nand (w_0624_, w_1096_, w_0082_);
xor (w_1114_, w_0302_, w_0461_);
xor (new_out5[0], w_0260_, w_0377_);
xor (w_1170_, w_1228_, w_0261_);
xor (w_0980_, w_0113_, w_0913_);
nor (new_out6[5], w_0964_, w_0314_);
nand (w_0540_, w_0397_, w_0586_);
and (w_0054_, w_0409_, w_0146_);
not (w_0717_, w_0588_);
nand (w_0523_, w_0575_, w_0294_);
nand (w_0882_, w_0206_, w_0823_);
nand (w_0919_, w_1011_, w_0004_);
nand (w_0177_, w_1116_, w_0486_);
or (w_1150_, w_0934_, w_0263_);
nand (w_0124_, w_0190_, w_0462_);
xor (w_0727_, new_in4[4], w_0317_);
xor (w_0930_, w_0469_, w_1031_);
or (w_0393_, new_out19[7], w_0489_);
xor (w_0027_, w_0987_, w_0264_);
nand (w_0921_, w_0361_, w_1114_);
nand (w_0312_, w_0399_, w_0655_);
nand (w_0654_, w_0986_, w_0565_);
xor (w_0105_, new_in6[4], w_0632_);
xor (new_out1[1], w_0619_, w_0562_);
xor (w_0448_, w_0882_, w_0795_);
nand (w_0398_, w_0925_, w_0618_);
xor (w_0110_, w_0907_, w_0144_);
nand (w_0039_, w_1071_, w_0655_);
xor (w_1206_, new_in14[0], w_1194_);
xor (w_0470_, new_in11[3], w_0734_);
nand (w_0590_, w_0399_, w_0577_);
xor (w_0513_, new_in5[2], w_0270_);
or (w_1073_, w_0027_, w_0347_);
nand (new_out3[2], w_0580_, w_0897_);
nand (w_1047_, w_0116_, w_0032_);
nand (w_1076_, w_1028_, w_0104_);
nand (w_0591_, w_0076_, w_0120_);
nand (w_0091_, w_0333_, w_0184_);
nand (w_0735_, w_0302_, w_0461_);
xor (w_0093_, new_in2[2], w_0037_);
nand (w_1130_, w_0028_, w_0262_);
xor (new_out7[5], w_0194_, w_0204_);
xor (new_out9[7], w_0884_, w_0466_);
xor (new_out16[5], w_0694_, w_0207_);
nand (w_0972_, new_in15[6], w_0354_);
and (w_0807_, w_0658_, w_0648_);
xor (w_0251_, new_in12[1], w_0909_);
xor (w_0837_, w_0821_, w_0160_);
xor (w_0063_, new_in9[2], w_0159_);
nand (w_0944_, w_0578_, w_0089_);
and (w_0155_, w_0584_, w_0229_);
nand (new_out3[0], w_1140_, w_0221_);
and (w_0551_, w_0950_, w_0322_);
xor (w_1220_, w_1017_, w_0045_);
xor (w_0305_, w_1063_, w_0161_);
xor (w_0883_, new_in15[6], w_0354_);
xor (w_0508_, w_1173_, w_0740_);
nand (w_1098_, w_0962_, w_0535_);
and (w_0342_, new_in2[0], w_0650_);
xor (w_0739_, w_0040_, w_0328_);
nand (w_0360_, w_0785_, w_0623_);
and (w_0387_, w_0725_, w_1002_);
xor (w_0218_, w_0858_, w_0054_);
nand (w_0171_, w_0096_, w_0420_);
nand (w_0664_, w_0538_, w_0848_);
nand (w_0353_, new_in14[2], w_0768_);
xor (w_1222_, w_0030_, w_1018_);
not (w_0634_, w_0422_);
xor (w_1171_, w_0355_, w_0073_);
not (new_out13[6], w_0303_);
and (w_0170_, w_0205_, w_0707_);
xor (w_0771_, w_1096_, w_0082_);
xor (w_0694_, w_0188_, w_0230_);
or (new_out15[6], w_0987_, w_0721_);
nand (w_0114_, new_in9[3], w_0671_);
nand (w_1131_, w_0447_, w_0296_);
nand (w_0520_, w_0837_, w_1100_);
xor (w_1044_, new_in1[5], w_0480_);
xor (new_out18[1], w_0436_, w_1128_);
xor (w_0585_, w_0721_, w_0029_);
nand (new_out24[6], w_0357_, w_0910_);
xor (w_0325_, w_0774_, w_1114_);
not (w_0269_, w_0848_);
xor (w_0244_, new_in11[4], w_0839_);
nand (w_0130_, w_0318_, w_0530_);
xor (w_1133_, w_0401_, w_0012_);
nand (w_1228_, w_0972_, w_0510_);
or (w_1116_, w_0168_, w_0059_);
xor (new_out9[0], w_0490_, w_0479_);
nand (w_0982_, w_0946_, w_0614_);
xor (new_out22[4], w_1167_, w_0566_);
nand (w_0647_, new_in12[2], w_0384_);
or (w_0025_, w_0696_, w_0422_);
xor (w_0282_, w_1084_, w_0256_);
xor (w_0289_, w_0356_, w_0407_);
xor (new_out14[3], w_0785_, w_0031_);
nand (w_0534_, w_0371_, w_0898_);
xor (w_0344_, w_0809_, w_0379_);
nand (new_out3[1], w_0907_, w_1154_);
nand (w_0744_, w_0529_, w_1111_);
nand (w_0810_, new_in4[3], w_0959_);
nand (w_0635_, w_1192_, w_0831_);
xor (w_0707_, w_0548_, w_0871_);
xor (w_0328_, w_0889_, w_0987_);
nand (w_0699_, new_in10[2], w_0771_);
nand (w_0140_, w_0599_, w_0049_);
xor (new_out4[1], w_0305_, w_0020_);
xor (w_0285_, w_0927_, w_0207_);
or (w_0099_, w_0020_, w_0837_);
xor (new_out4[4], w_0079_, w_0431_);
nand (w_1102_, w_0630_, w_0072_);
xor (w_0550_, new_in1[1], w_1056_);
xor (w_1132_, w_0787_, w_1060_);
nand (w_0816_, w_1210_, w_0956_);
nand (w_0127_, w_1180_, w_0616_);
and (w_0226_, w_0920_, w_0956_);
and (w_0696_, w_0253_, w_0335_);
not (w_0712_, new_in4[4]);
nand (w_0340_, w_0776_, w_1146_);
xor (new_out22[2], w_0605_, w_1190_);
not (w_0858_, w_0895_);
and (new_out17[1], w_0500_, w_0399_);
nand (w_0047_, w_0192_, w_0534_);
and (w_0765_, w_0627_, w_0968_);
xor (new_out8[2], w_0325_, w_0974_);
nand (w_0925_, w_1224_, w_0681_);
xor (w_0769_, new_in11[0], w_0521_);
nand (w_1042_, w_0693_, w_0540_);
xor (w_0314_, w_1118_, w_0663_);
not (w_0045_, w_0674_);
xor (w_0186_, w_0272_, w_0825_);
xor (w_0049_, w_1084_, w_0517_);
or (w_0818_, w_0013_, w_0958_);
xor (w_0137_, w_1133_, w_1200_);
or (w_0046_, w_0188_, w_0602_);
nand (w_0397_, w_1196_, w_0541_);
nand (w_1122_, w_0121_, w_0928_);
xor (w_0942_, new_in2[5], w_0326_);
nand (w_0452_, w_0679_, w_1179_);
nand (new_out2[0], w_0805_, w_0318_);
xor (w_1161_, w_0116_, w_0993_);
nand (w_0345_, w_0305_, w_0606_);
not (w_0774_, w_0361_);
nand (w_1162_, new_in15[5], w_0748_);
and (w_0113_, new_in12[0], w_0223_);
nand (w_0064_, w_0716_, w_0050_);
xor (w_1015_, w_0186_, w_0592_);
not (w_0954_, w_0697_);
xor (w_0897_, w_0538_, w_0848_);
xor (new_out14[1], w_1128_, w_0430_);
nand (w_0644_, w_0637_, w_0519_);
xor (w_1140_, w_0852_, w_1148_);
or (w_0522_, new_in8[3], new_in7[3]);
nand (w_0392_, w_1202_, w_0254_);
xor (w_0538_, w_0361_, w_1114_);
nand (w_0822_, new_in5[7], w_0364_);
nand (w_0068_, w_0574_, w_0799_);
nand (w_1121_, w_0143_, w_0314_);
xor (w_0101_, new_in11[1], w_1083_);
nand (w_0817_, w_0431_, w_0467_);
nand (w_1007_, w_1221_, w_0217_);
xor (new_out20[3], w_0380_, w_0442_);
nand (w_0050_, w_0311_, w_0576_);
nand (w_0992_, w_0783_, w_1189_);
and (w_0309_, new_out23[0], w_0429_);
xor (w_0210_, w_0006_, w_0414_);
xor (w_0596_, new_in14[3], w_0337_);
nor (w_0948_, w_0696_, w_1182_);
xor (w_0180_, w_0141_, w_0436_);
or (w_0372_, w_0425_, w_1220_);
xor (w_0401_, new_in10[1], w_0048_);
xor (w_0077_, new_in10[1], w_0669_);
xor (new_out5[2], w_0139_, w_0875_);
nand (w_0703_, w_0805_, w_0103_);
xor (w_0224_, w_0131_, w_0926_);
xor (w_1185_, w_0064_, w_0274_);
nand (w_0378_, new_in15[7], w_0943_);
or (w_0200_, w_0690_, w_0629_);
xor (w_0317_, w_1039_, w_0105_);
nand (w_0484_, w_0114_, w_1003_);
nand (w_0166_, w_0113_, w_0913_);
xor (w_0204_, w_1105_, w_0927_);
xor (w_0700_, w_0766_, w_0926_);
xor (w_0988_, w_0172_, w_0896_);
not (w_0673_, w_0426_);
nand (w_0182_, w_0058_, w_1088_);
and (w_0230_, w_0602_, w_0886_);
nand (w_0103_, w_0318_, w_0442_);
nand (w_0862_, w_0339_, w_0786_);
nor (w_0806_, w_0720_, w_1147_);
nand (w_0169_, w_0515_, w_0797_);
xor (new_out11[4], w_0754_, w_0931_);
xor (w_0141_, w_0505_, w_0755_);
nand (w_0976_, w_0902_, w_0864_);
nand (w_0653_, w_0092_, w_0572_);
xor (w_0704_, w_0869_, w_1032_);
nand (w_1088_, w_1098_, w_1101_);
nand (w_0636_, w_0056_, w_0392_);
xor (new_out1[0], w_0246_, w_0490_);
xor (w_0268_, new_in3[2], new_in16[2]);
xor (w_0724_, w_0620_, w_0580_);
xor (w_0768_, w_0477_, w_0410_);
nand (w_0545_, w_0626_, w_1109_);
xor (w_0697_, w_0683_, w_0162_);
nand (w_0098_, w_0987_, w_0456_);
xor (new_out4[0], w_0907_, w_0152_);
xor (w_0072_, new_in12[5], w_1062_);
xor (w_0681_, w_0332_, w_1126_);
or (w_0936_, w_1034_, w_0557_);
nand (w_0315_, w_1144_, w_1153_);
nand (w_0213_, new_in9[6], w_1080_);
and (w_0347_, w_0741_, w_1005_);
nand (w_0151_, new_in2[5], w_0326_);
nand (w_0831_, w_0485_, w_0242_);
nand (w_0267_, w_0610_, w_1125_);
xor (w_0661_, w_0177_, w_0224_);
or (w_1101_, w_1118_, w_1140_);
xor (w_0678_, w_0526_, w_0997_);
and (w_0813_, w_0750_, w_0008_);
nand (w_1163_, w_0889_, w_0987_);
xor (w_0788_, w_0290_, w_0044_);
nand (w_0183_, new_in6[3], w_0460_);
xor (w_0899_, w_1202_, w_0254_);
nand (w_0686_, w_0233_, w_0938_);
or (w_0612_, w_0876_, w_0595_);
nand (w_0090_, w_0798_, w_0708_);
xor (w_0865_, w_1079_, w_0468_);
xor (w_0277_, new_in13[4], w_0778_);
nand (w_0709_, w_0436_, w_1071_);
xor (new_out1[5], w_1191_, w_0285_);
nand (w_0938_, w_0833_, w_0483_);
nand (w_0043_, w_0785_, w_0301_);
nand (w_0973_, w_0484_, w_0308_);
xor (w_1030_, w_0186_, w_0449_);
xor (new_out18[4], w_0907_, w_0678_);
nand (w_0153_, w_0020_, w_0623_);
and (w_1013_, w_0453_, w_0432_);
xor (new_out10[3], w_0491_, w_0279_);
xor (new_out21[0], w_0388_, w_0202_);
nand (w_1127_, w_0042_, w_0077_);
or (w_0772_, w_0895_, w_0054_);
nand (w_0150_, w_0528_, w_0561_);
nand (w_0454_, w_1204_, w_0818_);
nand (w_0866_, w_0863_, w_0095_);
nand (w_1072_, w_0512_, w_0324_);
nand (w_1075_, new_in10[1], w_0669_);
xor (w_0115_, w_0068_, w_1213_);
and (w_0501_, w_0582_, w_1055_);
nand (w_0741_, w_0305_, w_1105_);
not (w_0355_, new_in11[5]);
nand (w_1111_, w_1072_, w_0257_);
xor (new_out22[6], w_0940_, w_0585_);
nand (w_0764_, w_0623_, w_0399_);
nand (w_1079_, w_1054_, w_0316_);
nand (w_1077_, w_0882_, w_0795_);
xor (w_0041_, w_1084_, w_0857_);
and (w_0915_, w_1163_, w_0236_);
nand (w_0844_, w_1136_, w_0446_);
and (w_0604_, w_0693_, w_0586_);
xor (w_0274_, w_1224_, w_1141_);
or (w_0283_, w_0186_, w_0449_);
xor (w_0620_, w_0607_, w_0216_);
nand (w_0902_, w_0822_, w_0516_);
nand (w_0334_, w_0728_, w_0265_);
and (w_0719_, w_0227_, w_0812_);
xor (w_0002_, new_in4[3], w_0959_);
not (w_0494_, w_0530_);
xor (new_out4[3], w_0857_, w_1105_);
nand (w_0782_, w_0869_, w_1032_);
nand (w_0292_, w_1128_, w_1205_);
nand (w_1050_, w_0940_, w_0585_);
xor (w_0273_, new_in2[5], w_0682_);
xor (new_out2[3], w_1174_, w_0944_);
not (w_0264_, w_0431_);
and (new_out17[3], w_0207_, w_1205_);
and (new_out17[2], w_0246_, w_0178_);
nand (w_0173_, w_0811_, w_0848_);
xor (new_out19[7], w_0857_, w_1224_);
nand (w_1117_, w_0754_, w_0931_);
xor (w_0333_, w_0399_, w_0577_);
nand (w_0376_, w_0353_, w_0009_);
nand (w_0477_, w_1075_, w_1127_);
nand (w_1191_, w_0283_, w_0088_);
xor (w_1154_, w_0436_, w_1071_);
or (w_0674_, w_1008_, w_0719_);
nand (w_0941_, new_in15[3], w_1143_);
nand (w_0720_, w_0143_, w_0807_);
xor (w_1165_, w_0592_, w_1230_);
nand (w_0614_, w_1001_, w_0727_);
nand (w_0679_, new_in5[4], w_0704_);
xor (w_0820_, new_in8[1], new_in7[1]);
nand (w_0779_, w_0649_, w_0636_);
xor (w_0029_, w_0637_, w_0519_);
and (w_1124_, w_1169_, w_0911_);
nand (w_0081_, w_0469_, w_1031_);
or (w_0579_, w_0852_, w_1148_);
nand (w_0362_, w_0982_, w_1175_);
xor (w_0038_, w_0250_, w_0445_);
nand (w_0846_, w_0995_, w_0646_);
nand (w_0640_, w_0070_, w_0549_);
nand (w_1106_, new_in2[4], w_0556_);
nand (w_0368_, w_0178_, w_0592_);
or (w_1055_, new_in16[7], new_in3[7]);
xor (w_0116_, w_1147_, w_0245_);
xor (w_0310_, new_in5[5], w_0189_);
xor (w_0216_, w_0197_, w_1123_);
nand (w_0809_, w_0286_, w_0854_);
nand (w_0983_, new_in6[2], w_0788_);
xor (w_0424_, w_0027_, w_0347_);
xor (new_out13[3], w_0837_, w_0927_);
nand (w_0975_, w_1151_, w_0352_);
xor (new_out22[0], w_0707_, w_0770_);
nand (w_1210_, w_0176_, w_0846_);
xor (w_1018_, new_in2[3], w_0790_);
xor (w_0352_, w_0785_, w_0301_);
nand (w_0176_, new_in13[2], w_0684_);
xor (w_0319_, w_0814_, w_1035_);
or (w_0805_, w_0079_, w_0422_);
and (w_0335_, w_0196_, w_0067_);
xor (w_1183_, w_0304_, w_0875_);
xor (w_0949_, new_in16[6], new_in3[2]);
xor (new_out23[5], new_out13[2], w_0955_);
nand (w_0761_, w_0655_, w_0701_);
not (w_1009_, w_0718_);
nand (w_0887_, new_in9[7], w_0369_);
xor (w_0399_, w_1000_, w_0935_);
nand (w_1129_, w_0343_, w_0428_);
nand (w_0657_, w_0872_, w_0093_);
not (w_0131_, w_1084_);
nand (w_0350_, w_1084_, w_0517_);
nand (w_0516_, w_1226_, w_0855_);
xor (w_0852_, w_0717_, w_0989_);
and (w_0833_, w_0207_, w_0500_);
xor (w_1126_, w_1013_, w_1199_);
xor (w_0449_, w_0634_, w_1220_);
nand (w_1176_, w_0172_, w_0896_);
xor (w_1027_, new_in15[1], w_0794_);
xor (new_out9[2], w_0190_, w_0462_);
xor (w_0785_, w_0525_, w_0212_);
xor (w_0663_, w_0630_, w_0072_);
nand (w_1107_, w_0052_, w_0698_);
and (w_0617_, w_0761_, w_0010_);
nand (w_1166_, w_0775_, w_1224_);
nand (w_0214_, new_in13[7], w_0154_);
nand (w_0728_, w_0659_, w_1142_);
nand (w_0389_, w_0787_, w_1060_);
nand (w_0543_, w_0923_, w_0295_);
nand (w_1104_, w_1140_, w_0021_);
xor (w_0524_, new_in2[6], w_0722_);
xor (w_0928_, new_in9[5], w_0403_);
or (w_0071_, w_0208_, w_0583_);
xor (w_0526_, w_0811_, w_0269_);
xor (w_0729_, new_in10[5], w_0413_);
xor (w_0730_, new_in11[3], w_0174_);
nand (new_out3[5], w_0500_, w_1134_);
nand (w_1003_, w_1034_, w_0557_);
xor (w_0128_, w_0872_, w_0093_);
nand (w_0109_, w_0552_, w_0238_);
nand (w_0860_, new_in14[5], w_0645_);
nand (w_1040_, w_0817_, w_0455_);
or (w_1177_, w_0987_, w_0264_);
or (w_0412_, w_0076_, w_0939_);
nand (w_0557_, w_0815_, w_1217_);
xor (w_0628_, new_in5[1], w_0705_);
xor (new_out4[5], w_0038_, w_1224_);
xor (w_0037_, w_0881_, w_0268_);
nand (w_0847_, w_1048_, w_0686_);
and (w_1120_, new_out2[0], w_0367_);
and (w_0052_, new_in11[0], w_0521_);
xor (w_0301_, w_1120_, w_1172_);
nand (w_0605_, w_0043_, w_0975_);
nand (w_1046_, w_1081_, w_0715_);
nand (w_0318_, w_0079_, w_0422_);
xor (w_0304_, w_0116_, w_0331_);
nand (w_1202_, w_0609_, w_0167_);
xor (w_0106_, w_0592_, w_0752_);
xor (w_1036_, w_0837_, w_1100_);
xor (w_0968_, w_1169_, w_0911_);
xor (w_0468_, new_in10[4], w_0001_);
and (new_out6[7], w_1224_, w_0606_);
nand (w_0965_, w_1036_, w_0929_);
xor (new_out2[2], w_0829_, w_0423_);
xor (w_1113_, w_0954_, w_0108_);
xor (w_0904_, w_0907_, w_0229_);
xor (w_0688_, w_0730_, w_0932_);
xor (w_0242_, new_in1[4], w_0676_);
nand (w_1226_, w_0784_, w_0826_);
xor (w_0684_, w_0300_, w_0834_);
xor (w_0384_, w_0728_, w_0265_);
xor (w_0521_, new_in8[0], new_in7[0]);
nand (w_0146_, w_1147_, w_0229_);
and (w_0191_, w_0132_, w_0209_);
xor (w_0296_, new_in16[5], new_in3[5]);
and (w_0835_, w_0039_, w_1146_);
nand (w_0118_, new_in11[5], w_0073_);
xor (w_1083_, new_in8[2], new_in7[1]);
xor (w_0763_, w_0371_, w_0898_);
nand (w_1019_, new_in2[6], w_0722_);
xor (w_0438_, w_0085_, w_0907_);
nand (w_0937_, new_in11[4], w_0839_);
xor (w_0488_, w_0580_, w_0163_);
and (w_0994_, new_in14[0], w_1194_);
or (w_0893_, w_0476_, w_0164_);
xor (w_0560_, new_in9[3], new_in13[3]);
xor (w_0229_, w_0642_, w_0467_);
nand (w_0804_, w_0605_, w_1190_);
not (w_0964_, w_1105_);
nand (w_0288_, w_1164_, w_0135_);
xor (w_0748_, w_0452_, w_0310_);
nand (w_0280_, new_in12[5], w_1062_);
xor (w_0957_, new_in1[7], w_1170_);
or (new_out15[2], w_0538_, w_0678_);
xor (new_out9[4], w_0181_, w_0906_);
nand (w_0033_, w_0491_, w_0279_);
or (new_out15[5], w_0305_, w_0615_);
xor (w_0655_, w_0987_, w_0673_);
xor (new_out11[0], w_1140_, w_0431_);
and (new_out17[4], w_0074_, w_0367_);
not (w_1211_, w_0875_);
xor (w_0074_, w_0677_, w_0739_);
xor (new_out9[1], w_1070_, w_0563_);
xor (w_0583_, w_1133_, w_0449_);
nand (w_0510_, w_0711_, w_0883_);
nand (w_0766_, w_0598_, w_0406_);
nand (w_0643_, w_0026_, w_0209_);
xor (new_out21[3], w_1104_, w_0381_);
xor (w_0517_, new_in15[6], new_in1[6]);
nand (w_0627_, w_0291_, w_0195_);
or (w_0552_, w_0314_, w_0218_);
xor (w_0207_, w_0454_, w_0668_);
nand (w_0385_, new_in14[3], w_0337_);
xor (w_0714_, w_0042_, w_0077_);
nor (new_out6[2], w_0974_, w_0449_);
nand (new_out24[4], w_1094_, w_0767_);
xor (w_0829_, w_1037_, w_0848_);
xor (w_0723_, new_in10[3], w_0149_);
xor (w_0337_, w_0842_, w_0471_);
xor (w_0432_, w_0627_, w_0968_);
xor (w_0354_, w_1076_, w_0239_);
xor (w_0931_, w_0848_, w_0592_);
xor (w_1095_, w_1072_, w_0257_);
or (w_0421_, w_0537_, w_0951_);
nand (w_0009_, w_0290_, w_0044_);
xor (w_1071_, new_in11[5], w_0141_);
or (w_0010_, w_0655_, w_0701_);
or (w_1214_, w_0020_, w_0623_);
not (w_0126_, new_in4[2]);
xor (w_0500_, w_0079_, w_0020_);
xor (new_out10[7], w_0078_, w_1048_);
nand (w_1201_, w_0673_, w_1205_);
xor (w_0556_, w_1042_, w_1181_);
xor (w_0461_, new_in15[0], new_in1[0]);
xor (w_0562_, w_0780_, w_1205_);
xor (new_out24[3], new_out10[3], w_0075_);
nand (w_0241_, w_0829_, w_0793_);
and (w_0737_, w_0069_, w_1029_);
xor (w_0446_, w_0235_, w_0918_);
or (w_0089_, w_0829_, w_0423_);
xor (w_0303_, w_0245_, w_0721_);
not (w_0407_, w_0109_);
xor (w_0755_, new_in9[1], w_0555_);
xor (w_0917_, w_0205_, w_0707_);
xor (new_out24[7], new_out10[7], w_0661_);
xor (w_0410_, new_in10[2], w_0771_);
xor (w_0756_, new_in2[0], w_0650_);
xor (new_out16[0], w_0987_, w_0490_);
nand (w_0594_, w_0417_, w_0185_);
nand (w_0032_, w_0175_, w_0564_);
not (w_1182_, w_0560_);
nand (w_0652_, w_0620_, w_0580_);
nand (w_0005_, w_1052_, w_1055_);
nor (w_0584_, w_0173_, w_0314_);
xor (new_out24[5], new_out10[5], w_0218_);
nand (w_1068_, w_1155_, w_0038_);
and (w_1218_, w_0058_, w_1101_);
and (w_1167_, w_0520_, w_0965_);
xor (w_0308_, new_in9[4], w_1138_);
nand (w_0797_, w_0960_, w_1063_);
and (w_0083_, new_in4[0], w_0880_);
xor (w_0951_, w_1178_, w_0259_);
and (w_1000_, w_0591_, w_0299_);
xor (w_0913_, new_in12[1], w_0148_);
nand (w_0828_, w_0292_, w_0847_);
nand (w_0692_, w_0761_, w_0481_);
nand (w_1038_, w_0477_, w_0410_);
not (w_0188_, w_0307_);
nand (w_0512_, w_0907_, w_0144_);
xor (w_0800_, w_0992_, w_0981_);
nand (w_0321_, w_0907_, w_0780_);
and (w_1212_, w_0205_, w_0246_);
xor (new_out9[3], w_0333_, w_0184_);
and (w_0811_, w_1139_, w_1071_);
nand (w_1045_, w_0232_, w_0483_);
nand (w_0869_, w_0933_, w_0062_);
nand (w_1085_, w_0546_, w_0527_);
and (w_0619_, w_0246_, w_0490_);
xor (new_out24[1], w_0945_, new_out10[1]);
nand (w_0787_, w_0808_, w_0327_);
xor (w_0313_, w_0692_, w_1165_);
nand (w_0133_, w_0908_, w_0522_);
nand (w_1082_, w_0487_, w_1223_);
xor (w_0433_, w_0623_, w_0399_);
xor (w_0873_, w_0092_, w_0572_);
xor (w_0632_, w_0440_, w_0900_);
xor (w_0911_, w_1046_, w_0055_);
xor (w_0263_, w_0615_, w_0234_);
and (w_1137_, w_0606_, w_0155_);
xor (w_0211_, w_0450_, w_0411_);
nand (w_0197_, w_1087_, w_0905_);
or (w_0950_, w_0325_, w_0974_);
nand (w_0731_, w_0500_, w_1049_);
xor (new_out16[1], w_0857_, w_0780_);
xor (w_0682_, new_in3[1], new_in16[5]);
nand (w_0918_, w_0573_, w_0976_);
or (w_0586_, new_in16[3], new_in3[3]);
xor (w_0912_, new_in5[3], w_0802_);
nand (w_0095_, w_0117_, w_1027_);
nand (w_0306_, w_0300_, w_0834_);
xor (new_out9[6], w_0247_, w_0323_);
nand (w_0329_, new_in4[5], w_0800_);
xor (w_0144_, w_0672_, new_out8[1]);
nand (w_0996_, w_0848_, w_0592_);
xor (w_0615_, w_0542_, w_0532_);
and (new_out6[6], w_0431_, w_0229_);
xor (w_0759_, w_0841_, w_0856_);
xor (new_out2[4], w_0116_, w_0032_);
not (w_0814_, new_in11[4]);
xor (w_0221_, w_0841_, w_0422_);
and (new_out6[1], w_0623_, w_0673_);
xor (w_0706_, w_1155_, w_0251_);
xor (new_out20[2], new_out19[7], w_0489_);
nand (w_0240_, w_0084_, w_0779_);
xor (w_0875_, w_0269_, w_0926_);
nand (w_0631_, w_0588_, w_0989_);
nand (w_0474_, w_0920_, w_0816_);
xor (new_out11[5], w_1160_, w_0916_);
xor (w_0004_, new_in6[3], w_0460_);
and (w_1178_, w_0060_, w_0641_);
xor (w_0457_, new_in3[3], new_in16[7]);
xor (w_0431_, w_0723_, w_0513_);
nand (w_0803_, w_0670_, w_0458_);
nand (w_0276_, w_0280_, w_1102_);
nand (w_0515_, w_0642_, w_0463_);
nand (w_0429_, w_0368_, w_0742_);
xor (w_0966_, w_0876_, w_0595_);
nand (w_0575_, new_in1[6], w_1022_);
xor (new_out7[3], w_0587_, w_0990_);
xor (w_0365_, w_0503_, w_0963_);
nand (w_1065_, w_0131_, w_0857_);
xor (w_0366_, w_0205_, w_0987_);
xor (w_0544_, new_in4[1], w_0873_);
nand (w_0287_, w_0152_, w_0367_);
and (w_0359_, w_0496_, w_0099_);
xor (w_0272_, w_0137_, w_0020_);
not (w_0021_, w_0314_);
nand (w_0084_, new_in5[3], w_1222_);
nand (w_0018_, w_0342_, w_0597_);
xor (new_out2[1], w_0318_, w_0530_);
xor (w_0189_, w_0942_, w_0539_);
xor (w_0935_, w_1098_, w_1218_);
xor (w_0154_, w_0523_, w_0957_);
not (w_0507_, w_0076_);
or (w_0209_, new_in8[5], new_in7[5]);
xor (w_1128_, w_0508_, w_0492_);
nand (w_0278_, w_0907_, w_0229_);
nand (w_1087_, w_0879_, w_0436_);
xor (w_0749_, w_0453_, w_0432_);
nand (w_0531_, new_in13[6], w_0344_);
xor (w_0677_, w_1203_, w_0558_);
nand (w_0767_, new_out10[4], w_0304_);
xor (w_0462_, w_0620_, w_1095_);
and (w_0466_, w_0656_, w_0187_);
xor (w_0363_, w_0076_, w_1037_);
and (w_0536_, new_in1[0], w_0427_);
and (w_0672_, w_0710_, w_0205_);
nand (w_0026_, w_0035_, w_0594_);
nor (w_0338_, w_0592_, w_0528_);
nand (w_0955_, w_0360_, w_0129_);
nand (w_0656_, w_0074_, w_0211_);
or (new_out15[0], w_0710_, w_0707_);
nand (w_0791_, w_0193_, w_0978_);
and (w_0051_, new_in8[0], new_in7[0]);
xor (w_1100_, w_0690_, w_0629_);
nand (w_0165_, w_0122_, w_0571_);
xor (w_1198_, w_0857_, w_0673_);
xor (new_out12[4], w_1147_, w_0801_);
xor (w_0867_, new_in14[1], w_0714_);
nand (w_0638_, w_0582_, w_0005_);
xor (new_out18[0], w_0710_, w_0074_);
xor (w_0926_, new_in4[5], w_0868_);
xor (new_out8[5], w_0305_, w_1105_);
xor (new_out12[6], w_0349_, w_0266_);
xor (w_0367_, w_0143_, w_0264_);
xor (new_out16[3], w_0038_, w_0399_);
not (w_1197_, new_out8[3]);
xor (new_out9[5], w_0838_, w_0434_);
xor (w_0577_, w_0744_, w_0617_);
xor (w_0849_, w_0002_, w_1016_);
and (w_0076_, w_0733_, w_0781_);
nor (w_0554_, w_1140_, w_0020_);
nor (w_0381_, w_0837_, w_0655_);
nand (w_1069_, w_0694_, w_0021_);
or (w_0578_, w_1037_, w_0269_);
xor (w_1103_, new_out13[7], w_0661_);
nand (w_0582_, new_in16[7], new_in3[7]);
xor (w_0162_, new_in9[7], new_in13[7]);
not (w_0793_, w_0611_);
xor (w_0456_, w_0696_, w_0889_);
xor (w_0246_, w_0038_, w_1133_);
xor (w_1209_, w_0416_, w_0359_);
xor (w_0427_, new_in15[0], w_1092_);
xor (w_0270_, new_in2[6], w_0949_);
nand (w_0708_, w_0619_, w_0562_);
nand (w_0250_, w_0350_, w_0140_);
xor (new_out4[2], w_0987_, w_1133_);
not (w_0710_, w_0841_);
xor (w_0266_, w_0311_, w_0576_);
and (w_0505_, new_in9[0], w_0830_);
nand (w_1096_, w_0293_, w_1107_);
xor (w_0475_, w_0170_, w_0439_);
xor (new_out23[0], w_0207_, w_0500_);
xor (w_0123_, w_0220_, w_1103_);
xor (new_out23[1], w_0833_, w_0483_);
xor (w_0563_, w_0780_, w_0827_);
nand (w_1086_, new_in2[2], w_0037_);
nand (w_0122_, w_0569_, w_1006_);
xor (w_0827_, w_0198_, w_0110_);
nor (w_0732_, w_0246_, w_0721_);
nand (w_1025_, w_0068_, w_1213_);
xor (w_0075_, w_0877_, w_1174_);
xor (w_1225_, w_0889_, w_0094_);
nand (w_0815_, new_in9[2], w_0159_);
xor (new_out18[3], w_1140_, w_0785_);
xor (w_0160_, w_0173_, w_0314_);
nand (w_0851_, w_0721_, w_0029_);
and (w_0117_, new_in15[0], w_1092_);
xor (w_0607_, w_0507_, w_0874_);
xor (w_0963_, new_in6[2], w_0788_);
or (w_1093_, w_0758_, w_1161_);
nand (w_1026_, w_0536_, w_0550_);
nand (w_0908_, w_0136_, w_0165_);
nand (w_0502_, w_0252_, w_0374_);
xor (w_1224_, w_1207_, w_0912_);
nand (w_0529_, w_0580_, w_0901_);
nand (w_0206_, w_0785_, w_0673_);
nand (w_0142_, w_0436_, w_0673_);
xor (new_out16[4], w_1037_, w_0178_);
nand (w_1097_, w_0305_, w_0964_);
nand (w_1169_, w_0860_, w_1025_);
xor (w_0850_, w_0096_, w_0420_);
nand (w_0541_, w_0881_, w_0268_);
and (w_0059_, w_0772_, w_0372_);
xor (w_0572_, new_in6[1], w_1014_);
xor (w_0718_, w_0633_, w_0747_);
not (w_0228_, w_1139_);
and (w_0690_, w_0685_, w_0612_);
xor (w_1141_, w_0282_, w_0700_);
nand (w_0984_, new_in9[4], w_1138_);
xor (w_0265_, new_in4[2], w_0365_);
nand (w_1020_, w_1219_, w_0495_);
nor (w_1021_, w_1205_, w_1141_);
xor (w_0259_, w_1136_, w_0446_);
nand (w_1039_, w_0183_, w_0919_);
nor (w_1053_, w_0580_, w_0678_);
xor (new_out16[2], w_0079_, w_0620_);
nand (w_0587_, w_0287_, w_0127_);
and (w_1174_, w_0175_, w_1110_);
xor (w_0668_, w_1149_, w_0737_);
nand (w_1180_, w_1201_, w_0593_);
nand (w_0060_, w_0214_, w_0391_);
not (w_0889_, w_0930_);
xor (w_0139_, w_0639_, w_0584_);
xor (w_0839_, w_0417_, w_0185_);
xor (new_out20[4], w_0530_, w_0703_);
xor (w_0616_, w_0152_, w_0367_);
nand (w_0465_, w_0640_, w_0613_);
xor (w_0721_, w_0702_, w_0514_);
or (w_0409_, w_0116_, w_0331_);
xor (w_0780_, w_0111_, w_0179_);
nand (w_0035_, new_in8[4], new_in7[4]);
xor (w_0646_, new_in13[2], w_0684_);
nand (w_0609_, new_in5[1], w_0705_);
xor (w_0841_, w_0696_, w_0560_);
nand (w_0320_, w_0503_, w_0963_);
xor (w_0239_, new_in5[6], w_0011_);
xor (w_0580_, w_0205_, w_0305_);
and (w_0878_, w_0953_, w_0844_);
not (w_0598_, w_0349_);
xor (w_0734_, new_in8[4], new_in7[3]);
nor (w_0443_, w_0907_, w_0785_);
nand (w_0057_, w_0764_, w_0297_);
nand (w_0633_, w_0887_, w_0243_);
nand (w_0648_, w_0363_, w_0499_);
xor (w_0801_, w_0476_, w_0164_);
xor (w_0262_, w_0907_, w_0780_);
and (w_0476_, w_0496_, w_0792_);
nand (w_0187_, w_0247_, w_0323_);
xor (new_out18[2], w_0538_, w_0707_);
not (w_0152_, w_0974_);
xor (w_1060_, new_in15[3], w_1143_);
xor (new_out1[3], w_0433_, w_1041_);
xor (w_0369_, w_1215_, w_0601_);
nand (w_0070_, w_0907_, w_1224_);
nand (w_1024_, w_0321_, w_1130_);
xor (w_0073_, w_0026_, w_0191_);
nand (w_1016_, w_0112_, w_0334_);
xor (w_0107_, w_0829_, w_0611_);
nand (w_0910_, new_out10[6], w_0134_);
nand (w_0733_, w_0537_, w_0951_);
nand (w_1152_, w_0137_, w_0020_);
xor (new_out12[0], w_0079_, w_0917_);
xor (w_1172_, w_0623_, w_0034_);
and (w_0395_, w_0631_, w_0579_);
nand (w_0294_, w_0809_, w_0379_);
nand (w_0416_, w_0472_, w_1077_);
nand (w_1157_, w_1078_, w_0524_);
nand (w_0284_, w_1084_, w_0857_);
xor (w_0906_, w_0186_, w_0313_);
nand (w_0482_, new_in9[5], w_0403_);
nand (w_0203_, w_0304_, w_1211_);
xor (w_0383_, new_in9[7], w_0369_);
not (w_0665_, w_0927_);
xor (new_out10[1], w_0028_, w_0262_);
xor (w_1017_, new_in12[4], w_0493_);
nand (w_0175_, w_0143_, w_0021_);
and (w_0537_, w_0633_, w_0747_);
xor (w_1008_, new_in12[3], w_0662_);
nand (w_0112_, new_in4[2], w_0365_);
nor (new_out6[4], w_0758_, w_0875_);
nand (w_0125_, w_1105_, w_0615_);
xor (w_0205_, w_0718_, w_0248_);
xor (new_out8[0], w_0710_, w_0205_);
xor (w_0903_, new_in10[5], w_0319_);
xor (w_1115_, new_in3[1], new_in16[1]);
xor (w_0003_, new_out19[7], w_0375_);
xor (new_out13[1], w_0785_, w_0623_);
nand (w_0324_, w_0198_, w_0110_);
or (w_0299_, w_0076_, w_0874_);
xor (w_0989_, new_in1[1], new_in15[1]);
nand (w_0339_, w_1186_, w_1065_);
nand (w_0863_, new_in15[1], w_0794_);
nand (w_0447_, w_0330_, w_0504_);
nand (w_0888_, w_1105_, w_0663_);
xor (w_0108_, new_in15[2], new_in1[2]);
xor (w_1031_, new_in9[6], w_1080_);
and (new_out6[0], w_0205_, w_0367_);
or (w_0357_, new_out10[6], w_0134_);
buf (new_out19[5:0], new_out8);
buf (new_out20[0], new_out8[5]);
endmodule

module new_sub_module3(
    input wire [1:0] new_in1,
    input wire [1:0] new_in10,
    input wire [1:0] new_in11,
    input wire [1:0] new_in12,
    input wire [1:0] new_in13,
    input wire [1:0] new_in14,
    input wire [1:0] new_in15,
    input wire [1:0] new_in2,
    input wire [1:0] new_in3,
    input wire [1:0] new_in4,
    input wire [1:0] new_in5,
    input wire [1:0] new_in6,
    input wire [1:0] new_in7,
    input wire [1:0] new_in8,
    input wire [1:0] new_in9,
    output wire new_out1,
    output wire new_out10,
    output wire new_out11,
    output wire new_out12,
    output wire new_out13,
    output wire new_out14,
    output wire new_out15,
    output wire new_out2,
    output wire new_out3,
    output wire new_out4,
    output wire new_out5,
    output wire new_out6,
    output wire new_out7,
    output wire new_out8,
    output wire new_out9
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
wire w_060_;
wire w_061_;
wire w_062_;
wire w_063_;
wire w_064_;
wire w_065_;
wire w_066_;
wire w_067_;
wire w_068_;
wire w_069_;
wire w_070_;
wire w_071_;
wire w_072_;
wire w_073_;
wire w_074_;
wire w_075_;
wire w_076_;
wire w_077_;
wire w_078_;
wire w_079_;
wire w_080_;
wire w_081_;
wire w_082_;
wire w_083_;
wire w_084_;
wire w_085_;
wire w_086_;
wire w_087_;
wire w_088_;
wire w_089_;
wire w_090_;
wire w_091_;
wire w_092_;
wire w_093_;
wire w_094_;
wire w_095_;
wire w_096_;
wire w_097_;
wire w_098_;
wire w_099_;
wire w_100_;
wire w_101_;
wire w_102_;
wire w_103_;
wire w_104_;
wire w_105_;
wire w_106_;
wire w_107_;
wire w_108_;
wire w_109_;
wire w_110_;
wire w_111_;
wire w_112_;
wire w_113_;
wire w_114_;
wire w_115_;
wire w_116_;
wire w_117_;
wire w_118_;
wire w_119_;
wire w_120_;
wire w_121_;
wire w_122_;
wire w_123_;
wire w_124_;
wire w_125_;
wire w_126_;
wire w_127_;
wire w_128_;
wire w_129_;
wire w_130_;
wire w_131_;
wire w_132_;
wire w_133_;
wire w_134_;
wire w_135_;
wire w_136_;
wire w_137_;
wire w_138_;
wire w_139_;
wire w_140_;
wire w_141_;
wire w_142_;
wire w_143_;
wire w_144_;
wire w_145_;
wire w_146_;
wire w_147_;
wire w_148_;
wire w_149_;
wire w_150_;
wire w_151_;
wire w_152_;
wire w_153_;
wire w_154_;
wire w_155_;
wire w_156_;
wire w_157_;
wire w_158_;
wire w_159_;
wire w_160_;
wire w_161_;
wire w_162_;
wire w_163_;
wire w_164_;
wire w_165_;
wire w_166_;
wire w_167_;
wire w_168_;
wire w_169_;
wire w_170_;
wire w_171_;
wire w_172_;
wire w_173_;
wire w_174_;
wire w_175_;
wire w_176_;
wire w_177_;
xor (w_074_, w_007_, w_023_);
xor (w_169_, new_in7[0], w_115_);
xor (w_090_, w_108_, w_084_);
xor (w_031_, w_176_, w_102_);
xor (w_144_, w_010_, w_094_);
and (w_161_, new_in1[1], new_in14[0]);
and (w_069_, new_in10[0], new_in12[0]);
xor (w_087_, new_in7[0], w_058_);
xor (w_132_, w_122_, w_128_);
xor (w_112_, w_114_, w_028_);
xor (w_166_, w_162_, w_005_);
and (w_078_, new_in1[0], new_in14[0]);
nor (w_129_, new_in12[0], new_in10[1]);
xor (w_085_, new_in10[1], new_in12[1]);
xor (w_050_, w_134_, w_110_);
xor (new_out2, w_141_, w_020_);
or (w_113_, new_in8[1], new_in3[0]);
xor (w_038_, w_172_, w_052_);
xor (w_020_, new_in7[0], w_166_);
and (w_097_, new_in4[1], new_in2[0]);
xor (w_174_, w_177_, w_069_);
nand (w_168_, new_in3[1], new_in8[0]);
xor (w_128_, w_019_, w_101_);
xor (w_055_, new_in7[0], w_042_);
xor (w_071_, w_160_, w_135_);
xor (w_094_, w_171_, w_006_);
xor (w_116_, w_079_, w_013_);
or (w_003_, new_in2[1], new_in4[1]);
or (w_143_, new_in11[1], new_in6[0]);
xor (w_160_, w_043_, w_027_);
xor (w_057_, w_124_, w_120_);
and (w_146_, w_102_, w_070_);
or (w_124_, new_in1[0], new_in14[1]);
xor (w_119_, new_in11[0], new_in6[0]);
nor (w_033_, w_129_, w_072_);
xor (w_047_, w_145_, w_133_);
xor (w_064_, w_136_, w_149_);
xor (new_out11, w_141_, w_123_);
xor (w_040_, w_062_, w_035_);
xor (w_013_, w_137_, w_165_);
xor (w_022_, w_078_, w_017_);
xor (new_out8, w_141_, w_169_);
xor (w_026_, w_059_, w_011_);
nor (w_100_, new_in5[0], new_in9[1]);
xor (w_091_, w_099_, w_001_);
xor (w_061_, new_in7[0], w_015_);
xor (new_out7, w_141_, w_154_);
nor (w_134_, w_175_, w_044_);
xor (w_138_, w_167_, w_148_);
xor (w_163_, new_in11[1], new_in6[0]);
and (w_000_, new_in5[0], new_in9[1]);
xor (w_109_, w_079_, w_144_);
xor (w_017_, w_103_, w_038_);
nand (w_172_, new_in13[1], new_in15[0]);
xor (w_008_, w_096_, w_053_);
xor (w_011_, new_in1[1], new_in14[1]);
xor (w_030_, w_126_, new_in5[1]);
xor (w_009_, w_124_, w_109_);
xor (w_136_, w_104_, w_086_);
xor (w_173_, w_156_, w_025_);
xor (w_005_, w_167_, w_032_);
xor (w_002_, w_100_, w_139_);
or (w_170_, new_in9[0], new_in5[1]);
xor (w_077_, w_019_, w_022_);
xor (w_117_, new_in7[0], w_118_);
xor (w_046_, w_131_, w_176_);
xor (w_098_, w_163_, w_067_);
nor (w_073_, new_in8[1], new_in3[1]);
xor (w_148_, w_078_, w_012_);
xor (w_150_, w_074_, w_155_);
and (w_122_, new_in6[1], new_in11[1]);
xor (w_105_, w_089_, w_119_);
xor (w_037_, w_134_, w_077_);
or (w_043_, new_in4[0], new_in2[0]);
xor (new_out3, new_in7[1], w_087_);
xor (w_083_, new_in2[1], new_in4[1]);
xor (new_out1, w_141_, w_061_);
nor (w_156_, new_in15[1], new_in13[1]);
xor (w_154_, new_in7[0], w_132_);
and (w_167_, w_019_, w_089_);
or (w_056_, new_in1[1], new_in14[1]);
nor (w_106_, w_161_, w_145_);
xor (w_028_, w_073_, w_006_);
nor (w_080_, new_in15[1], new_in13[0]);
xor (w_004_, w_140_, w_051_);
xor (w_075_, new_in7[0], w_098_);
xor (w_121_, w_163_, w_150_);
xor (w_152_, new_in7[0], w_147_);
xor (w_032_, w_161_, w_116_);
xor (w_036_, w_096_, w_174_);
xor (new_out12, w_141_, w_065_);
xor (w_115_, w_041_, w_130_);
xor (w_058_, w_175_, w_138_);
xor (w_133_, w_043_, w_008_);
xor (w_151_, w_155_, w_076_);
xor (w_140_, w_095_, w_082_);
xor (w_153_, w_063_, w_039_);
not (w_126_, new_in9[0]);
nor (w_145_, new_in1[1], new_in14[0]);
xor (w_039_, new_in4[0], new_in2[0]);
nor (w_120_, w_100_, w_000_);
xor (w_155_, new_in9[0], new_in5[0]);
xor (w_096_, new_in15[1], new_in13[0]);
xor (w_035_, w_003_, w_048_);
nand (w_104_, new_in10[0], new_in12[1]);
xor (new_out14, w_141_, w_092_);
xor (w_059_, w_097_, w_142_);
xor (new_out6, w_141_, w_055_);
xor (w_034_, new_in13[0], new_in15[0]);
xor (w_158_, w_021_, w_151_);
or (w_088_, new_in3[1], new_in8[0]);
xor (w_147_, w_051_, w_014_);
xor (w_018_, new_in7[0], w_029_);
xor (w_025_, w_177_, w_033_);
xor (w_082_, w_164_, w_145_);
xor (new_out15, new_in7[1], w_117_);
not (w_141_, new_in7[1]);
or (w_131_, new_in10[1], new_in12[1]);
xor (new_out13, w_141_, w_081_);
or (w_102_, new_in10[0], new_in12[1]);
xor (w_068_, new_in7[0], w_158_);
xor (w_125_, w_155_, w_026_);
xor (w_076_, w_056_, w_091_);
xor (w_051_, new_in6[1], new_in11[1]);
xor (new_out10, w_141_, w_075_);
xor (new_out9, w_141_, w_068_);
or (w_137_, new_in13[1], new_in15[0]);
and (w_041_, new_in11[0], new_in6[0]);
not (w_049_, new_in1[0]);
xor (w_081_, new_in7[0], w_121_);
nor (w_107_, new_in10[0], new_in12[0]);
or (w_159_, new_in4[0], new_in2[1]);
xor (w_142_, w_146_, w_080_);
xor (w_007_, w_093_, w_046_);
xor (w_048_, w_034_, w_045_);
nor (w_006_, w_107_, w_069_);
xor (w_054_, new_in4[1], new_in2[0]);
xor (w_024_, w_153_, w_031_);
xor (w_053_, w_168_, w_085_);
and (w_070_, w_088_, w_104_);
xor (w_065_, new_in7[0], w_050_);
xor (w_110_, w_170_, w_127_);
nor (w_175_, new_in6[1], new_in11[0]);
or (w_162_, new_in11[0], new_in6[0]);
xor (w_027_, w_114_, w_157_);
xor (w_101_, w_111_, w_090_);
xor (w_123_, new_in7[0], w_037_);
or (w_019_, new_in5[1], new_in9[1]);
and (w_176_, w_088_, w_168_);
xor (w_103_, new_in4[0], new_in2[1]);
xor (w_029_, w_122_, w_002_);
xor (w_067_, w_040_, w_000_);
xor (w_139_, w_062_, w_024_);
xor (w_127_, w_011_, w_016_);
nand (w_089_, new_in5[1], new_in9[1]);
xor (w_042_, w_047_, w_105_);
xor (w_135_, w_161_, w_030_);
xor (w_012_, w_097_, w_112_);
xor (w_001_, w_034_, w_066_);
xor (w_108_, w_049_, new_in14[0]);
nor (w_010_, new_in13[1], new_in15[0]);
xor (w_111_, w_063_, w_083_);
xor (new_out4, new_in7[1], w_152_);
and (w_072_, new_in12[0], new_in10[1]);
xor (w_165_, w_129_, w_171_);
xor (w_062_, new_in1[0], new_in14[1]);
xor (w_016_, w_003_, w_036_);
nand (w_177_, new_in8[0], new_in3[0]);
xor (w_023_, w_159_, w_106_);
and (w_095_, new_in9[0], new_in5[1]);
nor (w_086_, w_073_, w_060_);
and (w_044_, new_in6[1], new_in11[0]);
xor (w_052_, w_113_, w_072_);
nand (w_063_, new_in15[1], new_in13[1]);
xor (w_084_, w_113_, w_107_);
xor (w_114_, new_in15[1], new_in13[1]);
xor (w_130_, w_064_, w_057_);
xor (w_157_, w_107_, w_060_);
xor (w_149_, w_137_, w_054_);
and (w_060_, new_in8[1], new_in3[1]);
and (w_099_, new_in4[0], new_in2[1]);
xor (w_118_, w_044_, w_071_);
xor (w_015_, w_143_, w_125_);
and (w_079_, new_in2[1], new_in4[1]);
nand (w_093_, new_in13[0], new_in15[0]);
xor (w_164_, w_103_, w_173_);
xor (w_045_, w_177_, w_131_);
and (w_021_, new_in11[1], new_in6[0]);
xor (w_014_, w_100_, w_009_);
xor (w_171_, new_in8[1], new_in3[0]);
xor (new_out5, new_in7[1], w_018_);
xor (w_092_, new_in7[0], w_004_);
xor (w_066_, w_177_, w_085_);
endmodule
