module top_module (
    input wire        in1_sub_module1,
    input wire        in2_sub_module1,
    input wire        in3_sub_module1,
    input wire        in4_sub_module1,
    input wire        in5_sub_module1,
    input wire        in6_sub_module1,
    input wire        in7_sub_module1,
    input wire        in8_sub_module1,
    input wire        in9_sub_module1,
    input wire        in10_sub_module1,
    input wire        in11_sub_module1,
    input wire        in12_sub_module1,
    input wire        in13_sub_module1,
    input wire        in14_sub_module1,
    input wire        in15_sub_module1,
    input wire        in16_sub_module1,
    output wire       out1_sub_module1,
    output wire       out2_sub_module1,
    output wire       out3_sub_module1,
    output wire       out4_sub_module1,
    output wire       out5_sub_module1,
    output wire       out6_sub_module1,
    output wire       out7_sub_module1,
    output wire       out8_sub_module1,
    output wire       out9_sub_module1,
    output wire       out10_sub_module1,
    input wire  [5:0] in1_sub_module2,
    input wire  [5:0] in2_sub_module2,
    input wire  [5:0] in3_sub_module2,
    input wire  [5:0] in4_sub_module2,
    input wire  [5:0] in5_sub_module2,
    input wire  [5:0] in6_sub_module2,
    input wire  [5:0] in7_sub_module2,
    input wire  [5:0] in8_sub_module2,
    input wire  [7:0] in9_sub_module2,
    input wire  [7:0] in10_sub_module2,
    input wire  [7:0] in11_sub_module2,
    input wire  [7:0] in12_sub_module2,
    input wire  [7:0] in13_sub_module2,
    input wire  [7:0] in14_sub_module2,
    input wire  [7:0] in15_sub_module2,
    input wire  [7:0] in16_sub_module2,
    output wire [5:0] out1_sub_module2,
    output wire [5:0] out2_sub_module2,
    output wire [5:0] out3_sub_module2,
    output wire [5:0] out4_sub_module2,
    output wire [5:0] out5_sub_module2,
    output wire [5:0] out6_sub_module2,
    output wire [5:0] out7_sub_module2,
    output wire [5:0] out8_sub_module2,
    output wire [5:0] out9_sub_module2,
    output wire [5:0] out10_sub_module2,
    output wire [5:0] out11_sub_module2,
    output wire [5:0] out12_sub_module2,
    output wire [7:0] out13_sub_module2,
    output wire [7:0] out14_sub_module2,
    output wire [7:0] out15_sub_module2,
    output wire [7:0] out16_sub_module2,
    output wire [7:0] out17_sub_module2,
    output wire [7:0] out18_sub_module2,
    output wire [7:0] out19_sub_module2,
    output wire [7:0] out20_sub_module2,
    output wire [7:0] out21_sub_module2,
    output wire [7:0] out22_sub_module2,
    output wire [7:0] out23_sub_module2,
    output wire [7:0] out24_sub_module2,
    input wire  [1:0] in1_sub_module3,
    input wire  [1:0] in2_sub_module3,
    input wire  [1:0] in3_sub_module3,
    input wire  [1:0] in4_sub_module3,
    input wire  [1:0] in5_sub_module3,
    input wire  [1:0] in6_sub_module3,
    input wire  [1:0] in7_sub_module3,
    input wire  [1:0] in8_sub_module3,
    input wire  [1:0] in9_sub_module3,
    input wire  [1:0] in10_sub_module3,
    input wire  [1:0] in11_sub_module3,
    input wire  [1:0] in12_sub_module3,
    input wire  [1:0] in13_sub_module3,
    input wire  [1:0] in14_sub_module3,
    input wire  [1:0] in15_sub_module3,
    output wire       out1_sub_module3,
    output wire       out2_sub_module3,
    output wire       out3_sub_module3,
    output wire       out4_sub_module3,
    output wire       out5_sub_module3,
    output wire       out6_sub_module3,
    output wire       out7_sub_module3,
    output wire       out8_sub_module3,
    output wire       out9_sub_module3,
    output wire       out10_sub_module3,
    output wire       out11_sub_module3,
    output wire       out12_sub_module3,
    output wire       out13_sub_module3,
    output wire       out14_sub_module3,
    output wire       out15_sub_module3
);
    sub_module1 U1 (
        .in1(in1_sub_module1),
        .in2(in2_sub_module1),
        .in3(in3_sub_module1),
        .in4(in4_sub_module1),
        .in5(in5_sub_module1),
        .in6(in6_sub_module1),
        .in7(in7_sub_module1),
        .in8(in8_sub_module1),
        .in9(in9_sub_module1),
        .in10(in10_sub_module1),
        .in11(in11_sub_module1),
        .in12(in12_sub_module1),
        .in13(in13_sub_module1),
        .in14(in14_sub_module1),
        .in15(in15_sub_module1),
        .in16(in16_sub_module1),
        .out1(out1_sub_module1),
        .out2(out2_sub_module1),
        .out3(out3_sub_module1),
        .out4(out4_sub_module1),
        .out5(out5_sub_module1),
        .out6(out6_sub_module1),
        .out7(out7_sub_module1),
        .out8(out8_sub_module1),
        .out9(out9_sub_module1),
        .out10(out10_sub_module1)
    );

    sub_module2 U2 (
        .in1(in1_sub_module2),
        .in2(in2_sub_module2),
        .in3(in3_sub_module2),
        .in4(in4_sub_module2),
        .in5(in5_sub_module2),
        .in6(in6_sub_module2),
        .in7(in7_sub_module2),
        .in8(in8_sub_module2),
        .in9(in9_sub_module2),
        .in10(in10_sub_module2),
        .in11(in11_sub_module2),
        .in12(in12_sub_module2),
        .in13(in13_sub_module2),
        .in14(in14_sub_module2),
        .in15(in15_sub_module2),
        .in16(in16_sub_module2),
        .out1(out1_sub_module2),
        .out2(out2_sub_module2),
        .out3(out3_sub_module2),
        .out4(out4_sub_module2),
        .out5(out5_sub_module2),
        .out6(out6_sub_module2),
        .out7(out7_sub_module2),
        .out8(out8_sub_module2),
        .out9(out9_sub_module2),
        .out10(out10_sub_module2),
        .out11(out11_sub_module2),
        .out12(out12_sub_module2),
        .out13(out13_sub_module2),
        .out14(out14_sub_module2),
        .out15(out15_sub_module2),
        .out16(out16_sub_module2),
        .out17(out17_sub_module2),
        .out18(out18_sub_module2),
        .out19(out19_sub_module2),
        .out20(out20_sub_module2),
        .out21(out21_sub_module2),
        .out22(out22_sub_module2),
        .out23(out23_sub_module2),
        .out24(out24_sub_module2)
    );

    sub_module3 U3 (
        .in1(in1_sub_module3),
        .in2(in2_sub_module3),
        .in3(in3_sub_module3),
        .in4(in4_sub_module3),
        .in5(in5_sub_module3),
        .in6(in6_sub_module3),
        .in7(in7_sub_module3),
        .in8(in8_sub_module3),
        .in9(in9_sub_module3),
        .in10(in10_sub_module3),
        .in11(in11_sub_module3),
        .in12(in12_sub_module3),
        .in13(in13_sub_module3),
        .in14(in14_sub_module3),
        .in15(in15_sub_module3),
        .out1(out1_sub_module3),
        .out2(out2_sub_module3),
        .out3(out3_sub_module3),
        .out4(out4_sub_module3),
        .out5(out5_sub_module3),
        .out6(out6_sub_module3),
        .out7(out7_sub_module3),
        .out8(out8_sub_module3),
        .out9(out9_sub_module3),
        .out10(out10_sub_module3),
        .out11(out11_sub_module3),
        .out12(out12_sub_module3),
        .out13(out13_sub_module3),
        .out14(out14_sub_module3),
        .out15(out15_sub_module3)
    );

endmodule
