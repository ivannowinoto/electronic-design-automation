module new_sub_module1(
    input wire [2:0] new_in1,
    input wire [2:0] new_in10,
    input wire [2:0] new_in12,
    input wire [2:0] new_in13,
    input wire [2:0] new_in2,
    input wire [2:0] new_in5,
    input wire [2:0] new_in7,
    input wire [3:0] new_in11,
    input wire [3:0] new_in14,
    input wire [3:0] new_in3,
    input wire [3:0] new_in4,
    input wire [3:0] new_in6,
    input wire [3:0] new_in8,
    input wire [3:0] new_in9,
    output wire [1:0] new_out10,
    output wire [1:0] new_out11,
    output wire [1:0] new_out3,
    output wire [1:0] new_out7,
    output wire [1:0] new_out9,
    output wire [2:0] new_out1,
    output wire [2:0] new_out2,
    output wire [2:0] new_out4,
    output wire [2:0] new_out5,
    output wire [2:0] new_out8,
    output wire [3:0] new_out12,
    output wire [3:0] new_out6
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
wire w_060_;
wire w_061_;
wire w_062_;
wire w_063_;
wire w_064_;
wire w_065_;
wire w_066_;
wire w_067_;
wire w_068_;
wire w_069_;
wire w_070_;
wire w_071_;
wire w_072_;
wire w_073_;
wire w_074_;
wire w_075_;
wire w_076_;
wire w_077_;
wire w_078_;
wire w_079_;
wire w_080_;
wire w_081_;
wire w_082_;
wire w_083_;
wire w_084_;
wire w_085_;
wire w_086_;
wire w_087_;
wire w_088_;
wire w_089_;
wire w_090_;
wire w_091_;
wire w_092_;
wire w_093_;
wire w_094_;
wire w_095_;
wire w_096_;
wire w_097_;
wire w_098_;
wire w_099_;
wire w_100_;
wire w_101_;
wire w_102_;
wire w_103_;
wire w_104_;
wire w_105_;
wire w_106_;
wire w_107_;
wire w_108_;
wire w_109_;
wire w_110_;
wire w_111_;
wire w_112_;
wire w_113_;
wire w_114_;
wire w_115_;
wire w_116_;
wire w_117_;
wire w_118_;
wire w_119_;
wire w_120_;
wire w_121_;
wire w_122_;
wire w_123_;
wire w_124_;
wire w_125_;
wire w_126_;
wire w_127_;
wire w_128_;
wire w_129_;
wire w_130_;
wire w_131_;
wire w_132_;
wire w_133_;
wire w_134_;
wire w_135_;
wire w_136_;
wire w_137_;
wire w_138_;
wire w_139_;
wire w_140_;
wire w_141_;
wire w_142_;
wire w_143_;
wire w_144_;
wire w_145_;
wire w_146_;
wire w_147_;
wire w_148_;
wire w_149_;
wire w_150_;
wire w_151_;
wire w_152_;
wire w_153_;
wire w_154_;
wire w_155_;
wire w_156_;
wire w_157_;
wire w_158_;
wire w_159_;
wire w_160_;
wire w_161_;
wire w_162_;
wire w_163_;
wire w_164_;
wire w_165_;
wire w_166_;
wire w_167_;
wire w_168_;
wire w_169_;
wire w_170_;
wire w_171_;
wire w_172_;
wire w_173_;
wire w_174_;
wire w_175_;
wire w_176_;
wire w_177_;
wire w_178_;
wire w_179_;
wire w_180_;
wire w_181_;
wire w_182_;
wire w_183_;
wire w_184_;
wire w_185_;
wire w_186_;
wire w_187_;
wire w_188_;
wire w_189_;
wire w_190_;
wire w_191_;
wire w_192_;
wire w_193_;
wire w_194_;
wire w_195_;
wire w_196_;
wire w_197_;
wire w_198_;
wire w_199_;
wire w_200_;
wire w_201_;
wire w_202_;
wire w_203_;
wire w_204_;
wire w_205_;
wire w_206_;
wire w_207_;
wire w_208_;
wire w_209_;
wire w_210_;
wire w_211_;
wire w_212_;
wire w_213_;
wire w_214_;
wire w_215_;
wire w_216_;
wire w_217_;
wire w_218_;
wire w_219_;
wire w_220_;
wire w_221_;
wire w_222_;
wire w_223_;
wire w_224_;
wire w_225_;
wire w_226_;
wire w_227_;
wire w_228_;
wire w_229_;
wire w_230_;
wire w_231_;
wire w_232_;
wire w_233_;
wire w_234_;
wire w_235_;
wire w_236_;
wire w_237_;
wire w_238_;
wire w_239_;
wire w_240_;
wire w_241_;
wire w_242_;
wire w_243_;
wire w_244_;
wire w_245_;
wire w_246_;
wire w_247_;
wire w_248_;
wire w_249_;
wire w_250_;
wire w_251_;
wire w_252_;
wire w_253_;
wire w_254_;
wire w_255_;
wire w_256_;
wire w_257_;
wire w_258_;
wire w_259_;
wire w_260_;
wire w_261_;
wire w_262_;
wire w_263_;
wire w_264_;
wire w_265_;
wire w_266_;
wire w_267_;
wire w_268_;
wire w_269_;
wire w_270_;
wire w_271_;
wire w_272_;
wire w_273_;
wire w_274_;
wire w_275_;
wire w_276_;
wire w_277_;
wire w_278_;
wire w_279_;
wire w_280_;
wire w_281_;
wire w_282_;
wire w_283_;
wire w_284_;
wire w_285_;
wire w_286_;
wire w_287_;
wire w_288_;
wire w_289_;
wire w_290_;
wire w_291_;
wire w_292_;
wire w_293_;
wire w_294_;
wire w_295_;
wire w_296_;
wire w_297_;
wire w_298_;
wire w_299_;
wire w_300_;
wire w_301_;
wire w_302_;
wire w_303_;
wire w_304_;
wire w_305_;
wire w_306_;
xor (w_077_, w_256_, w_181_);
xor (w_122_, new_in12[2], w_075_);
and (w_157_, w_251_, w_030_);
nand (w_144_, w_156_, w_250_);
xor (w_199_, new_in8[2], w_294_);
xor (w_131_, new_in9[0], new_in6[0]);
nand (w_031_, w_033_, w_238_);
and (w_212_, w_158_, w_047_);
xor (w_209_, w_147_, w_162_);
xor (new_out3[0], w_240_, w_208_);
xor (new_out12[2], w_084_, w_097_);
xor (w_105_, new_in14[1], w_139_);
and (w_271_, w_136_, w_073_);
xor (new_out11[0], w_109_, w_035_);
nand (w_081_, w_295_, w_082_);
xor (w_202_, w_175_, w_165_);
nand (w_088_, w_086_, w_232_);
xor (w_126_, new_in2[2], w_017_);
nand (w_001_, w_174_, w_044_);
nand (w_050_, w_265_, w_257_);
and (w_096_, w_207_, w_224_);
nand (w_044_, w_248_, w_199_);
xor (new_out2[2], w_009_, w_214_);
nand (w_221_, w_165_, w_054_);
xor (new_out10[0], w_143_, w_298_);
not (w_178_, w_243_);
xor (w_003_, new_in7[2], new_in10[2]);
nand (w_283_, w_125_, w_048_);
xor (w_161_, w_291_, w_254_);
xor (w_075_, w_260_, w_201_);
and (new_out5[1], w_088_, w_277_);
nand (w_037_, new_in9[3], new_in6[3]);
xor (w_189_, w_273_, w_245_);
nand (w_305_, w_200_, w_038_);
xor (new_out11[1], w_239_, w_000_);
and (new_out5[2], w_217_, w_286_);
xor (w_114_, w_127_, w_182_);
nand (w_036_, w_252_, w_144_);
not (w_193_, w_109_);
xor (w_195_, w_006_, w_187_);
xor (w_303_, w_060_, w_126_);
xor (w_112_, w_083_, w_205_);
xor (w_026_, w_092_, w_102_);
nand (w_200_, new_in4[1], new_in3[1]);
xor (w_151_, new_in4[1], new_in3[1]);
xor (w_268_, w_059_, w_281_);
xor (w_165_, w_172_, w_105_);
xor (w_008_, w_113_, w_104_);
xor (w_227_, new_in8[0], w_170_);
nand (w_021_, w_115_, w_133_);
nand (w_295_, w_274_, w_011_);
nand (w_028_, w_092_, w_163_);
xor (w_296_, w_285_, w_128_);
xor (new_out8[0], w_109_, w_208_);
xor (w_016_, w_295_, w_082_);
xor (new_out7[1], w_063_, w_293_);
xor (w_027_, new_in8[1], w_204_);
nand (w_207_, new_in1[1], w_261_);
nand (w_260_, w_107_, w_176_);
nand (w_060_, w_152_, w_020_);
xor (w_201_, new_in5[2], w_070_);
nand (w_238_, w_153_, w_228_);
xor (w_203_, new_in1[2], w_009_);
nand (w_002_, w_043_, w_109_);
nand (w_225_, w_103_, w_079_);
xor (w_236_, w_217_, w_286_);
xor (w_280_, w_248_, w_199_);
or (w_141_, w_096_, w_203_);
nand (w_150_, new_in1[2], w_114_);
nand (w_048_, w_010_, w_160_);
nand (w_072_, w_202_, w_240_);
xor (w_217_, w_056_, w_068_);
xor (w_233_, w_129_, w_045_);
or (w_242_, new_in1[1], w_261_);
xor (w_181_, new_in5[1], w_093_);
and (w_265_, w_189_, w_067_);
xor (w_245_, w_246_, w_145_);
xor (w_070_, w_196_, w_065_);
and (w_010_, new_in12[0], w_049_);
not (w_259_, w_127_);
nand (w_270_, w_072_, w_050_);
nand (w_138_, w_117_, w_306_);
and (w_121_, w_111_, w_237_);
nand (w_147_, w_087_, w_091_);
nand (w_158_, w_202_, w_003_);
xor (w_140_, w_180_, w_046_);
xor (w_043_, w_220_, w_264_);
xor (w_257_, w_202_, w_240_);
nand (new_out4[2], w_214_, w_121_);
nand (w_232_, w_080_, w_231_);
and (w_172_, new_in14[0], w_131_);
xor (w_041_, w_194_, w_173_);
xor (w_177_, new_in10[0], new_in1[0]);
nand (w_258_, new_in5[2], w_070_);
xor (w_206_, new_in4[2], new_in3[2]);
nand (w_005_, w_211_, w_124_);
xor (w_097_, w_161_, w_215_);
not (w_129_, w_275_);
not (w_123_, new_in1[0]);
xor (w_254_, new_in1[1], w_303_);
xor (w_046_, w_165_, w_054_);
xor (w_263_, new_in14[2], w_209_);
not (w_188_, w_233_);
nand (w_246_, w_262_, w_034_);
nand (w_069_, w_127_, w_303_);
xor (w_022_, new_in9[1], new_in6[1]);
nand (w_018_, w_113_, w_104_);
xor (w_162_, new_in6[2], new_in9[2]);
nand (w_134_, new_in2[2], w_017_);
nand (w_176_, w_256_, w_181_);
xor (w_017_, w_283_, w_122_);
xor (new_out6[1], w_190_, w_143_);
nand (w_107_, new_in5[1], w_093_);
nand (w_055_, w_161_, w_215_);
xor (w_067_, new_in9[0], new_in11[2]);
nor (w_063_, w_051_, w_013_);
nand (w_247_, w_101_, w_304_);
or (w_234_, w_156_, w_250_);
nand (w_211_, w_008_, w_041_);
nand (w_226_, w_221_, w_130_);
xor (w_143_, w_264_, w_182_);
xor (w_231_, w_003_, w_009_);
xor (w_065_, new_in1[2], new_in10[2]);
nand (w_120_, w_031_, w_269_);
nand (w_103_, new_in8[3], w_016_);
xor (w_304_, new_in10[1], new_in1[1]);
nand (w_169_, w_148_, w_081_);
nand (w_187_, w_258_, w_108_);
and (w_014_, new_in9[0], new_in6[0]);
xor (w_009_, w_259_, w_182_);
nand (w_108_, w_260_, w_201_);
nand (w_153_, w_025_, w_018_);
and (w_276_, w_055_, w_074_);
xor (w_013_, w_270_, w_218_);
nand (w_148_, new_in4[3], new_in3[3]);
xor (w_090_, w_251_, w_030_);
nand (w_095_, w_289_, w_089_);
xor (w_145_, w_169_, w_225_);
xor (w_064_, w_268_, w_296_);
nand (w_146_, w_275_, w_045_);
xor (w_298_, w_273_, w_116_);
nand (w_038_, w_272_, w_151_);
nand (new_out4[0], w_071_, w_051_);
xor (w_085_, new_in11[1], w_110_);
xor (w_035_, w_189_, w_067_);
xor (w_297_, w_026_, w_061_);
xor (w_049_, new_in5[0], w_177_);
xor (w_054_, w_230_, w_085_);
xor (w_015_, w_244_, w_029_);
xor (w_273_, new_in14[0], w_131_);
nand (w_174_, new_in8[2], w_294_);
nand (w_154_, new_in11[1], w_110_);
or (w_039_, w_026_, w_061_);
xor (w_082_, new_in4[3], new_in3[3]);
nand (w_047_, w_243_, w_137_);
nand (w_118_, w_302_, w_249_);
nand (w_255_, new_in10[1], new_in1[1]);
xor (w_099_, w_021_, w_271_);
nand (w_125_, new_in12[1], w_077_);
xor (new_out6[2], w_024_, w_112_);
xor (w_205_, w_008_, w_041_);
nand (w_224_, w_095_, w_242_);
xor (w_058_, new_in1[0], w_285_);
xor (w_269_, w_115_, w_133_);
xor (new_out1[0], new_in1[0], w_114_);
nand (w_124_, w_083_, w_205_);
xor (w_220_, w_278_, w_263_);
xor (w_299_, w_132_, w_166_);
xor (w_253_, w_092_, w_163_);
nand (w_155_, w_288_, w_078_);
nand (w_191_, w_155_, w_300_);
xor (new_out12[0], w_088_, w_277_);
nand (w_197_, new_in14[3], w_299_);
xor (w_109_, new_in10[0], new_in7[0]);
and (w_083_, w_264_, w_182_);
and (w_061_, w_002_, w_229_);
and (w_076_, w_028_, w_290_);
nand (w_237_, w_036_, w_222_);
xor (w_294_, w_305_, w_206_);
nand (w_079_, w_001_, w_284_);
xor (w_106_, w_005_, w_267_);
nand (w_056_, w_066_, w_086_);
xor (w_164_, w_010_, w_160_);
and (w_186_, w_207_, w_242_);
xor (new_out12[3], w_064_, w_276_);
nand (w_159_, w_005_, w_267_);
and (w_012_, w_193_, w_143_);
xor (w_170_, new_in4[0], new_in3[0]);
nand (w_292_, w_132_, w_166_);
nand (w_115_, w_134_, w_282_);
xor (w_094_, w_178_, w_137_);
xor (w_284_, new_in8[3], w_016_);
xor (w_228_, new_in7[2], new_in13[2]);
nand (w_252_, w_245_, w_090_);
xor (new_out2[0], w_043_, w_106_);
xor (new_out8[2], w_076_, w_149_);
nand (w_156_, w_198_, w_023_);
nand (w_053_, new_in12[2], w_075_);
and (w_080_, w_235_, w_039_);
and (w_167_, new_out5[1], w_236_);
xor (w_216_, w_036_, w_222_);
xor (w_062_, w_220_, w_015_);
xor (w_139_, w_014_, w_022_);
xor (w_004_, w_092_, w_112_);
nand (w_042_, w_057_, w_223_);
xor (new_out1[1], new_in1[1], w_285_);
and (w_272_, new_in4[0], new_in3[0]);
and (w_135_, new_in8[0], w_170_);
xor (w_183_, w_118_, w_098_);
xor (w_166_, new_in9[3], new_in6[3]);
nand (w_030_, w_197_, w_191_);
nand (w_007_, w_196_, w_065_);
xor (w_215_, w_096_, w_203_);
xor (w_277_, w_212_, w_168_);
nand (w_152_, new_in2[1], w_164_);
xor (w_092_, new_in10[1], new_in7[1]);
nand (w_251_, w_037_, w_292_);
nand (w_066_, w_003_, w_114_);
xor (new_out10[1], w_140_, w_112_);
nand (w_287_, w_172_, w_105_);
xor (w_149_, w_003_, w_071_);
xor (w_240_, new_in9[1], new_in11[3]);
nand (w_229_, w_270_, w_218_);
nand (w_100_, new_in8[1], w_204_);
nand (w_136_, w_006_, w_187_);
xor (w_261_, w_008_, w_185_);
nand (w_266_, w_283_, w_122_);
xor (new_out6[3], w_071_, w_106_);
xor (w_110_, w_135_, w_027_);
and (w_019_, w_120_, w_146_);
not (w_051_, w_106_);
nand (w_011_, w_305_, w_206_);
nand (w_006_, w_241_, w_007_);
nand (w_275_, w_069_, w_159_);
nand (w_020_, w_194_, w_173_);
xor (new_out12[1], new_out5[1], w_236_);
nand (w_052_, w_053_, w_266_);
xor (w_285_, w_041_, w_031_);
nand (w_175_, w_192_, w_032_);
xor (w_301_, w_001_, w_284_);
nand (w_132_, w_171_, w_119_);
xor (w_160_, new_in12[1], w_077_);
xor (w_133_, w_052_, w_195_);
xor (w_168_, w_123_, w_043_);
nand (w_032_, w_246_, w_145_);
xor (w_208_, w_226_, w_062_);
and (w_256_, new_in5[0], w_177_);
nand (w_171_, new_in6[2], new_in9[2]);
nand (w_196_, w_255_, w_247_);
xor (new_out1[2], new_in1[2], w_303_);
xor (w_267_, w_127_, w_303_);
and (w_291_, w_117_, w_306_);
nand (w_290_, w_142_, w_253_);
xor (w_173_, new_in2[1], w_164_);
nand (w_244_, w_154_, w_213_);
nand (w_025_, new_in7[1], new_in13[1]);
xor (new_out9[1], w_012_, w_004_);
nand (w_034_, w_118_, w_098_);
and (w_059_, w_179_, w_184_);
nand (w_117_, new_in1[0], w_285_);
xor (w_137_, w_202_, w_003_);
nand (w_288_, new_in14[2], w_209_);
nand (w_033_, new_in7[2], new_in13[2]);
and (w_101_, new_in10[0], new_in1[0]);
nand (w_306_, w_056_, w_058_);
nand (w_073_, w_052_, w_195_);
xor (w_029_, new_in11[2], w_280_);
xor (w_300_, new_in14[3], w_299_);
nand (w_078_, w_278_, w_263_);
xor (w_116_, new_in11[0], w_227_);
xor (w_098_, new_in11[3], w_301_);
and (w_142_, w_109_, w_208_);
nand (w_192_, w_169_, w_225_);
and (w_113_, new_in13[0], new_in7[0]);
nand (w_023_, w_042_, w_040_);
or (new_out4[1], w_188_, w_216_);
xor (w_093_, w_101_, w_304_);
and (w_180_, w_273_, w_116_);
xor (w_214_, w_099_, w_019_);
nand (w_074_, w_084_, w_097_);
and (w_128_, w_150_, w_141_);
and (w_243_, w_092_, w_189_);
xor (w_293_, w_233_, w_297_);
nand (w_213_, w_230_, w_085_);
xor (new_out7[0], w_051_, w_013_);
or (w_086_, w_080_, w_231_);
nand (w_111_, w_175_, w_157_);
nand (w_289_, new_in1[0], w_043_);
nand (w_223_, w_226_, w_062_);
not (w_068_, w_058_);
not (new_out6[0], w_140_);
nor (new_out5[0], w_297_, w_094_);
nand (w_274_, new_in4[2], new_in3[2]);
xor (w_127_, w_153_, w_228_);
nand (w_130_, w_180_, w_046_);
xor (new_out9[0], w_109_, w_143_);
xor (w_163_, w_042_, w_040_);
xor (w_222_, w_175_, w_157_);
and (w_194_, new_in2[0], w_219_);
xor (w_000_, w_265_, w_257_);
nand (w_184_, w_138_, w_254_);
and (w_230_, new_in11[0], w_227_);
xor (w_286_, w_095_, w_186_);
nand (w_087_, new_in9[1], new_in6[1]);
xor (w_239_, w_092_, w_189_);
nand (w_057_, w_220_, w_015_);
nand (w_210_, w_135_, w_027_);
xor (w_219_, new_in12[0], w_049_);
nand (w_282_, w_060_, w_126_);
xor (w_104_, new_in7[1], new_in13[1]);
nand (w_071_, w_144_, w_234_);
nand (w_119_, w_147_, w_162_);
xor (new_out3[1], w_109_, w_163_);
xor (new_out2[1], w_102_, w_233_);
xor (w_045_, w_031_, w_269_);
xor (w_218_, w_043_, w_109_);
nand (w_278_, w_279_, w_287_);
or (w_084_, new_out5[2], w_167_);
nand (w_241_, new_in1[2], new_in10[2]);
xor (w_182_, new_in2[0], w_219_);
nand (w_179_, new_in1[1], w_303_);
xor (w_250_, w_245_, w_090_);
nand (w_249_, w_244_, w_029_);
nand (w_279_, new_in14[1], w_139_);
nand (w_248_, w_100_, w_210_);
xor (w_264_, new_in13[0], new_in7[0]);
nand (w_302_, new_in11[2], w_280_);
nand (w_198_, w_185_, w_183_);
xor (w_185_, w_155_, w_300_);
xor (new_out8[1], w_142_, w_253_);
xor (w_204_, w_272_, w_151_);
not (w_190_, w_208_);
not (w_102_, w_261_);
nand (w_091_, w_014_, w_022_);
nand (w_262_, new_in11[3], w_301_);
nand (w_235_, w_092_, w_261_);
xor (w_281_, new_in1[2], w_269_);
not (w_024_, w_163_);
or (w_089_, w_212_, w_168_);
xor (w_040_, w_185_, w_183_);
endmodule

module new_sub_module2(
    input wire [1:0] new_in10,
    input wire [1:0] new_in15,
    input wire [1:0] new_in2,
    input wire [1:0] new_in6,
    input wire [1:0] new_in7,
    input wire [1:0] new_in8,
    input wire [1:0] new_in9,
    input wire [4:0] new_in1,
    input wire [4:0] new_in11,
    input wire [4:0] new_in12,
    input wire [4:0] new_in13,
    input wire [4:0] new_in14,
    input wire [4:0] new_in3,
    input wire [4:0] new_in4,
    input wire [4:0] new_in5,
    output wire [1:0] new_out1,
    output wire [1:0] new_out10,
    output wire [1:0] new_out5,
    output wire [1:0] new_out6,
    output wire [1:0] new_out9,
    output wire [2:0] new_out11,
    output wire [2:0] new_out12,
    output wire [2:0] new_out13,
    output wire [2:0] new_out3,
    output wire [2:0] new_out8,
    output wire [3:0] new_out14,
    output wire [3:0] new_out2,
    output wire [3:0] new_out4,
    output wire [3:0] new_out7
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
wire w_060_;
wire w_061_;
wire w_062_;
wire w_063_;
wire w_064_;
wire w_065_;
wire w_066_;
wire w_067_;
wire w_068_;
wire w_069_;
wire w_070_;
wire w_071_;
wire w_072_;
wire w_073_;
wire w_074_;
wire w_075_;
wire w_076_;
wire w_077_;
wire w_078_;
wire w_079_;
wire w_080_;
wire w_081_;
wire w_082_;
wire w_083_;
wire w_084_;
wire w_085_;
wire w_086_;
wire w_087_;
wire w_088_;
wire w_089_;
wire w_090_;
wire w_091_;
wire w_092_;
wire w_093_;
wire w_094_;
wire w_095_;
wire w_096_;
wire w_097_;
wire w_098_;
wire w_099_;
wire w_100_;
wire w_101_;
wire w_102_;
wire w_103_;
wire w_104_;
wire w_105_;
wire w_106_;
wire w_107_;
wire w_108_;
wire w_109_;
wire w_110_;
wire w_111_;
wire w_112_;
wire w_113_;
wire w_114_;
wire w_115_;
wire w_116_;
wire w_117_;
wire w_118_;
wire w_119_;
wire w_120_;
wire w_121_;
wire w_122_;
wire w_123_;
wire w_124_;
wire w_125_;
wire w_126_;
wire w_127_;
wire w_128_;
wire w_129_;
wire w_130_;
wire w_131_;
wire w_132_;
wire w_133_;
wire w_134_;
wire w_135_;
wire w_136_;
wire w_137_;
wire w_138_;
wire w_139_;
wire w_140_;
wire w_141_;
wire w_142_;
wire w_143_;
wire w_144_;
wire w_145_;
wire w_146_;
wire w_147_;
wire w_148_;
wire w_149_;
wire w_150_;
wire w_151_;
wire w_152_;
wire w_153_;
wire w_154_;
wire w_155_;
wire w_156_;
wire w_157_;
wire w_158_;
wire w_159_;
wire w_160_;
wire w_161_;
wire w_162_;
wire w_163_;
wire w_164_;
wire w_165_;
wire w_166_;
wire w_167_;
wire w_168_;
wire w_169_;
wire w_170_;
wire w_171_;
wire w_172_;
wire w_173_;
wire w_174_;
wire w_175_;
wire w_176_;
wire w_177_;
wire w_178_;
wire w_179_;
wire w_180_;
wire w_181_;
wire w_182_;
wire w_183_;
wire w_184_;
wire w_185_;
wire w_186_;
wire w_187_;
wire w_188_;
wire w_189_;
wire w_190_;
wire w_191_;
wire w_192_;
wire w_193_;
wire w_194_;
wire w_195_;
wire w_196_;
wire w_197_;
wire w_198_;
wire w_199_;
wire w_200_;
wire w_201_;
wire w_202_;
wire w_203_;
wire w_204_;
wire w_205_;
wire w_206_;
wire w_207_;
wire w_208_;
wire w_209_;
wire w_210_;
wire w_211_;
wire w_212_;
wire w_213_;
wire w_214_;
wire w_215_;
wire w_216_;
wire w_217_;
wire w_218_;
wire w_219_;
wire w_220_;
wire w_221_;
wire w_222_;
wire w_223_;
wire w_224_;
wire w_225_;
wire w_226_;
wire w_227_;
wire w_228_;
wire w_229_;
wire w_230_;
wire w_231_;
wire w_232_;
wire w_233_;
wire w_234_;
wire w_235_;
wire w_236_;
wire w_237_;
wire w_238_;
wire w_239_;
wire w_240_;
wire w_241_;
wire w_242_;
wire w_243_;
wire w_244_;
wire w_245_;
wire w_246_;
wire w_247_;
wire w_248_;
wire w_249_;
wire w_250_;
wire w_251_;
wire w_252_;
wire w_253_;
wire w_254_;
wire w_255_;
wire w_256_;
wire w_257_;
wire w_258_;
wire w_259_;
wire w_260_;
wire w_261_;
wire w_262_;
wire w_263_;
wire w_264_;
wire w_265_;
wire w_266_;
wire w_267_;
wire w_268_;
wire w_269_;
wire w_270_;
wire w_271_;
wire w_272_;
wire w_273_;
wire w_274_;
wire w_275_;
wire w_276_;
wire w_277_;
wire w_278_;
wire w_279_;
wire w_280_;
wire w_281_;
wire w_282_;
wire w_283_;
wire w_284_;
wire w_285_;
wire w_286_;
wire w_287_;
wire w_288_;
wire w_289_;
wire w_290_;
wire w_291_;
wire w_292_;
wire w_293_;
wire w_294_;
wire w_295_;
wire w_296_;
wire w_297_;
wire w_298_;
wire w_299_;
wire w_300_;
wire w_301_;
wire w_302_;
wire w_303_;
wire w_304_;
wire w_305_;
wire w_306_;
wire w_307_;
wire w_308_;
wire w_309_;
wire w_310_;
wire w_311_;
wire w_312_;
wire w_313_;
wire w_314_;
wire w_315_;
wire w_316_;
wire w_317_;
wire w_318_;
wire w_319_;
wire w_320_;
wire w_321_;
wire w_322_;
wire w_323_;
wire w_324_;
nand (w_172_, w_305_, w_257_);
nand (w_035_, w_198_, w_312_);
xor (new_out7[1], new_in15[1], w_180_);
nand (w_275_, w_211_, w_159_);
nand (w_063_, w_051_, w_295_);
nand (w_008_, w_000_, w_169_);
or (w_065_, w_112_, w_028_);
xor (w_180_, w_207_, w_204_);
or (w_264_, w_017_, w_181_);
xor (new_out14[0], w_239_, w_071_);
xor (w_160_, w_260_, w_318_);
xor (new_out7[2], new_in7[0], w_223_);
xor (w_118_, w_051_, w_295_);
nand (w_282_, w_133_, w_287_);
xor (new_out2[3], w_174_, w_218_);
xor (w_293_, w_179_, w_248_);
nand (w_289_, w_177_, w_323_);
xor (w_019_, w_002_, w_053_);
or (w_027_, w_203_, w_059_);
xor (w_186_, w_081_, w_298_);
and (w_083_, w_038_, w_202_);
nand (w_009_, w_165_, w_167_);
xor (w_229_, new_in14[3], w_293_);
xor (w_169_, w_186_, w_017_);
xor (w_042_, new_in5[4], w_032_);
nand (w_140_, w_056_, w_217_);
not (w_151_, w_091_);
xor (w_101_, new_in11[1], w_231_);
nand (w_077_, w_156_, w_269_);
nand (w_049_, w_069_, w_276_);
xor (w_244_, new_in10[1], new_in6[1]);
nand (w_154_, w_149_, w_185_);
nand (w_316_, new_in4[3], new_in13[3]);
nand (w_106_, w_112_, w_028_);
nand (w_062_, new_in14[3], w_293_);
nand (w_188_, w_289_, w_029_);
xor (w_156_, w_153_, w_190_);
xor (w_003_, w_203_, w_059_);
and (w_000_, w_111_, w_061_);
and (w_090_, new_in12[0], new_in3[0]);
xor (w_001_, w_134_, w_244_);
xor (new_out12[0], w_038_, w_096_);
nand (w_306_, w_120_, w_155_);
nand (w_176_, w_016_, w_089_);
nand (w_040_, new_in12[4], new_in3[4]);
xor (w_080_, new_in8[0], w_324_);
and (w_173_, w_079_, w_188_);
nand (w_290_, w_232_, w_221_);
nand (w_310_, w_137_, w_086_);
xor (w_133_, new_in11[3], w_023_);
nor (w_240_, w_036_, w_299_);
xor (w_258_, w_317_, w_238_);
xor (w_070_, w_085_, w_097_);
xor (w_268_, w_307_, w_220_);
nand (w_205_, w_117_, w_233_);
nand (w_305_, new_in4[1], new_in13[1]);
xor (w_018_, new_in11[4], w_127_);
xor (w_081_, w_067_, w_030_);
and (w_174_, w_153_, w_190_);
nand (w_320_, w_307_, w_220_);
nand (w_084_, w_195_, w_164_);
xor (w_250_, w_069_, w_161_);
not (w_053_, w_037_);
xor (w_097_, new_in3[3], new_in12[3]);
xor (w_164_, w_252_, w_021_);
nand (w_177_, new_in1[4], w_197_);
nand (w_227_, w_122_, w_031_);
xor (w_091_, w_016_, w_089_);
xor (w_046_, new_in7[0], new_in15[0]);
xor (w_135_, w_111_, w_317_);
xor (w_128_, w_214_, w_072_);
xor (w_112_, w_300_, w_299_);
and (w_004_, new_in11[0], w_012_);
xor (new_out12[2], w_206_, w_119_);
xor (w_292_, new_in14[4], w_130_);
xor (w_114_, w_247_, w_193_);
xor (new_out6[0], w_038_, w_215_);
xor (w_086_, new_in4[4], new_in13[4]);
nand (w_256_, new_in2[1], w_100_);
nand (w_182_, w_090_, w_094_);
xor (w_238_, w_215_, w_202_);
nand (w_108_, new_in1[3], w_138_);
nand (w_271_, w_143_, w_272_);
nor (w_236_, w_195_, w_164_);
xor (new_out8[0], w_318_, w_118_);
xor (new_out8[2], w_195_, w_219_);
nand (w_045_, w_315_, w_224_);
nand (w_192_, w_179_, w_248_);
nand (w_322_, w_107_, w_196_);
xor (w_214_, w_157_, w_018_);
nand (w_107_, w_260_, w_318_);
and (w_117_, new_in14[0], w_273_);
xor (w_222_, w_237_, w_123_);
and (w_150_, new_in5[0], w_104_);
nand (w_139_, w_124_, w_020_);
and (w_010_, new_in7[0], new_in15[0]);
nand (w_011_, w_243_, w_238_);
xor (w_037_, w_000_, w_169_);
nand (w_015_, w_108_, w_152_);
nand (w_257_, w_237_, w_123_);
xor (w_145_, new_in5[2], w_319_);
xor (w_295_, w_186_, w_195_);
xor (w_279_, new_in10[0], new_in6[0]);
and (w_199_, w_219_, w_005_);
and (w_208_, w_017_, w_260_);
xor (w_076_, w_226_, w_025_);
xor (w_158_, w_117_, w_233_);
xor (new_out13[0], w_080_, w_019_);
nand (w_274_, new_in4[4], new_in13[4]);
xor (w_220_, new_in14[2], w_183_);
xor (w_130_, w_137_, w_086_);
nand (w_148_, w_033_, w_251_);
nand (w_201_, w_194_, w_182_);
xor (new_out13[2], w_114_, w_113_);
xor (w_304_, w_206_, w_303_);
nand (w_034_, w_214_, w_021_);
nand (w_036_, w_263_, w_164_);
xor (w_219_, w_099_, w_288_);
xor (new_out4[1], w_014_, w_213_);
xor (new_out3[0], w_038_, w_202_);
xor (w_260_, w_206_, w_114_);
nand (w_321_, w_103_, w_042_);
xor (new_out1[1], w_064_, w_092_);
xor (new_out10[0], w_053_, w_135_);
xor (new_out14[3], w_013_, w_102_);
xor (w_017_, w_252_, w_254_);
xor (w_313_, w_239_, w_081_);
xor (w_012_, new_in5[0], w_104_);
xor (w_249_, w_250_, w_303_);
nand (w_323_, w_015_, w_171_);
nand (w_198_, new_in1[1], w_158_);
xor (w_100_, w_010_, w_088_);
nand (w_039_, w_322_, w_258_);
xor (w_082_, new_in11[2], w_129_);
xor (w_298_, w_124_, w_020_);
nand (w_228_, new_in8[1], w_168_);
nand (w_263_, w_011_, w_109_);
xor (new_out11[0], w_215_, w_208_);
xor (w_113_, w_278_, w_128_);
xor (w_127_, w_103_, w_042_);
xor (w_038_, new_in1[0], w_285_);
xor (w_248_, new_in4[3], new_in13[3]);
nand (w_115_, new_in11[3], w_023_);
nand (w_267_, w_201_, w_261_);
and (w_144_, w_306_, w_049_);
not (w_302_, w_287_);
nand (w_232_, w_013_, w_202_);
not (w_206_, w_050_);
nand (w_047_, w_274_, w_310_);
xor (w_058_, w_036_, w_299_);
xor (new_out11[2], w_156_, w_131_);
xor (w_031_, new_in9[1], w_001_);
xor (w_088_, new_in7[1], new_in15[1]);
xor (new_out2[2], w_211_, w_159_);
xor (w_273_, new_in4[0], new_in13[0]);
xor (w_014_, w_263_, w_164_);
nand (w_028_, w_084_, w_284_);
nand (w_187_, w_172_, w_286_);
and (w_051_, w_111_, w_317_);
nand (w_157_, w_115_, w_282_);
xor (w_129_, w_045_, w_145_);
xor (w_300_, w_250_, w_013_);
xor (w_147_, w_269_, w_266_);
xor (new_out2[1], w_280_, w_126_);
nand (w_216_, w_162_, w_320_);
xor (w_123_, new_in4[1], new_in13[1]);
xor (w_171_, new_in1[4], w_197_);
xor (w_212_, new_in12[4], new_in3[4]);
and (w_102_, w_058_, w_147_);
xor (new_out7[3], new_in7[1], w_230_);
nand (w_005_, w_284_, w_301_);
xor (w_023_, w_056_, w_217_);
xor (w_247_, w_234_, w_294_);
and (w_048_, w_002_, w_053_);
nand (w_152_, w_175_, w_148_);
nand (w_110_, new_in4[2], new_in13[2]);
xor (new_out4[0], w_219_, w_236_);
xor (w_074_, new_in1[2], w_268_);
nand (w_235_, new_in5[4], w_032_);
nand (w_315_, new_in5[1], w_314_);
xor (w_072_, w_322_, w_258_);
nand (w_218_, w_077_, w_275_);
nand (w_178_, w_245_, w_008_);
not (w_064_, w_318_);
xor (w_286_, new_in4[2], new_in13[2]);
nand (w_211_, w_044_, w_060_);
nand (w_242_, new_in10[1], new_in6[1]);
nand (w_055_, new_in5[3], w_070_);
and (w_006_, w_238_, w_318_);
or (w_078_, w_300_, w_299_);
nand (w_155_, w_235_, w_321_);
and (w_124_, new_in8[0], w_324_);
not (w_043_, w_156_);
xor (w_002_, w_121_, w_082_);
xor (w_276_, w_120_, w_155_);
nand (w_153_, w_066_, w_262_);
and (w_266_, w_078_, w_106_);
and (w_234_, w_242_, w_209_);
nand (w_085_, w_253_, w_267_);
xor (new_out9[1], new_in8[1], w_125_);
nand (w_116_, w_048_, w_003_);
nand (w_226_, w_151_, w_007_);
nand (w_170_, w_239_, w_081_);
not (w_189_, w_260_);
nand (w_026_, w_290_, w_270_);
or (w_301_, w_200_, w_283_);
xor (w_050_, w_035_, w_074_);
not (w_013_, w_203_);
xor (w_020_, new_in8[1], w_168_);
nand (w_283_, w_054_, w_039_);
xor (w_243_, w_141_, w_144_);
or (w_087_, w_300_, w_189_);
xor (w_223_, w_290_, w_270_);
not (w_141_, w_214_);
xor (w_119_, w_009_, w_309_);
and (w_134_, new_in10[0], new_in6[0]);
nand (w_167_, w_226_, w_025_);
and (w_105_, w_002_, w_238_);
xor (new_out3[1], w_083_, w_041_);
nand (w_022_, w_004_, w_101_);
xor (w_089_, w_300_, w_189_);
xor (w_297_, w_002_, w_050_);
xor (w_202_, w_175_, w_148_);
nand (w_125_, w_064_, w_072_);
nand (w_098_, new_in9[1], w_001_);
nand (w_073_, new_in11[1], w_231_);
and (w_142_, w_311_, w_052_);
nor (w_071_, w_151_, w_072_);
xor (w_285_, new_in14[0], w_273_);
xor (w_168_, w_122_, w_031_);
xor (w_075_, w_254_, w_050_);
nand (w_044_, w_252_, w_112_);
nand (w_272_, w_225_, w_292_);
nand (w_165_, w_037_, w_219_);
and (w_213_, w_300_, w_299_);
xor (w_255_, new_in5[1], w_314_);
and (w_122_, new_in9[0], w_279_);
and (w_193_, w_228_, w_139_);
nand (w_079_, w_047_, w_271_);
and (w_067_, new_in1[0], w_285_);
nand (w_068_, w_216_, w_229_);
xor (w_309_, w_014_, w_181_);
xor (new_out5[1], w_298_, w_105_);
xor (w_183_, w_172_, w_286_);
nand (w_225_, w_062_, w_068_);
and (w_095_, w_034_, w_026_);
xor (w_025_, w_037_, w_219_);
xor (w_303_, w_289_, w_029_);
and (w_149_, new_in2[0], w_046_);
nand (w_190_, w_256_, w_154_);
nand (w_146_, new_in14[1], w_222_);
xor (w_159_, w_156_, w_269_);
xor (w_217_, new_in5[3], w_070_);
nand (w_057_, w_163_, w_212_);
nand (w_287_, w_246_, w_259_);
nand (w_307_, w_146_, w_205_);
xor (w_175_, new_in1[3], w_138_);
xor (w_299_, w_043_, w_303_);
nand (w_296_, w_081_, w_021_);
xor (w_197_, w_225_, w_292_);
xor (new_out7[0], new_in15[0], w_297_);
xor (w_200_, w_195_, w_164_);
xor (w_288_, w_243_, w_238_);
xor (w_324_, new_in9[0], w_279_);
nand (w_191_, w_186_, w_195_);
and (w_131_, w_317_, w_164_);
nand (w_281_, w_085_, w_097_);
xor (new_out11[1], w_252_, w_006_);
xor (w_252_, w_149_, w_185_);
nand (w_056_, w_024_, w_166_);
xor (w_041_, w_081_, w_021_);
nand (w_137_, w_316_, w_192_);
xor (w_111_, w_080_, w_038_);
nand (w_278_, w_027_, w_116_);
xor (w_007_, w_111_, w_093_);
nand (w_109_, w_099_, w_288_);
not (w_161_, w_276_);
xor (w_231_, w_150_, w_255_);
xor (w_061_, w_215_, w_239_);
and (w_184_, w_014_, w_277_);
nand (w_265_, new_in11[4], w_127_);
xor (w_029_, w_047_, w_271_);
nand (w_060_, w_280_, w_126_);
nand (w_291_, w_157_, w_018_);
xor (w_230_, w_095_, w_249_);
nand (w_054_, w_317_, w_238_);
xor (w_185_, new_in2[1], w_100_);
nand (w_162_, new_in14[2], w_183_);
not (w_093_, w_061_);
nand (w_312_, w_067_, w_030_);
xor (w_021_, w_015_, w_171_);
xor (new_out10[1], w_181_, w_118_);
nand (w_099_, w_087_, w_176_);
and (w_294_, w_098_, w_227_);
xor (w_314_, w_090_, w_094_);
nand (w_262_, w_010_, w_088_);
nand (w_308_, new_in3[3], new_in12[3]);
nand (w_196_, w_178_, w_160_);
xor (w_270_, w_214_, w_021_);
nand (w_245_, w_186_, w_017_);
nand (w_209_, w_134_, w_244_);
xor (w_138_, w_216_, w_229_);
xor (w_318_, w_002_, w_156_);
and (w_132_, w_254_, w_260_);
nand (w_166_, w_045_, w_145_);
nand (w_246_, new_in11[2], w_129_);
nand (w_120_, w_040_, w_057_);
xor (w_311_, w_214_, w_144_);
xor (new_out13[1], w_298_, w_210_);
not (w_181_, w_059_);
nand (w_016_, w_191_, w_063_);
xor (new_out2[0], w_215_, w_200_);
nand (w_259_, w_121_, w_082_);
nand (w_121_, w_073_, w_022_);
xor (w_059_, w_178_, w_160_);
xor (w_233_, new_in14[1], w_222_);
xor (w_269_, w_311_, w_052_);
nand (w_179_, w_110_, w_187_);
xor (new_out3[2], w_136_, w_304_);
or (w_221_, w_207_, w_204_);
nand (w_103_, w_055_, w_140_);
nand (w_207_, w_002_, w_050_);
xor (w_204_, w_203_, w_202_);
xor (w_126_, w_252_, w_112_);
nand (w_069_, w_265_, w_291_);
and (w_237_, new_in4[0], new_in13[0]);
xor (w_203_, w_133_, w_302_);
xor (w_195_, w_002_, w_214_);
nand (w_241_, w_083_, w_041_);
xor (w_254_, w_004_, w_101_);
xor (new_out4[3], w_052_, w_240_);
nand (w_253_, new_in12[2], new_in3[2]);
xor (new_out8[1], w_317_, w_091_);
xor (new_out14[1], w_254_, w_199_);
nand (w_033_, new_in1[2], w_268_);
xor (w_030_, new_in1[1], w_158_);
xor (new_out4[2], w_142_, w_058_);
and (w_136_, w_296_, w_241_);
nand (w_194_, new_in12[1], new_in3[1]);
xor (w_317_, w_254_, w_013_);
xor (new_out12[1], w_081_, w_076_);
nand (w_277_, w_106_, w_065_);
xor (w_094_, new_in12[1], new_in3[1]);
nand (w_143_, new_in14[4], w_130_);
xor (w_096_, w_091_, w_007_);
xor (w_215_, new_in2[0], w_046_);
xor (new_out5[0], w_080_, w_132_);
xor (w_032_, w_163_, w_212_);
nand (w_251_, w_035_, w_074_);
and (w_280_, w_215_, w_200_);
xor (w_092_, w_170_, w_075_);
xor (w_052_, w_174_, w_173_);
nand (w_284_, w_200_, w_283_);
xor (new_out9[0], new_in8[0], w_264_);
xor (new_out14[2], w_002_, w_184_);
xor (new_out1[0], w_017_, w_313_);
xor (w_239_, new_in11[0], w_012_);
nand (w_224_, w_150_, w_255_);
xor (w_261_, new_in12[2], new_in3[2]);
xor (w_210_, w_048_, w_003_);
nand (w_066_, new_in7[1], new_in15[1]);
xor (new_out6[1], w_081_, w_252_);
nand (w_163_, w_308_, w_281_);
nand (w_024_, new_in5[2], w_319_);
xor (w_319_, w_201_, w_261_);
xor (w_104_, new_in12[0], new_in3[0]);
endmodule

module new_sub_module3(
    input wire [2:0] new_in3,
    input wire [2:0] new_in6,
    input wire [2:0] new_in8,
    input wire [3:0] new_in4,
    input wire [3:0] new_in5,
    input wire [3:0] new_in7,
    input wire [4:0] new_in1,
    input wire [4:0] new_in12,
    input wire [4:0] new_in9,
    input wire [5:0] new_in11,
    input wire [5:0] new_in15,
    input wire [5:0] new_in2,
    input wire [6:0] new_in10,
    input wire [6:0] new_in13,
    input wire [6:0] new_in14,
    output wire [1:0] new_out1,
    output wire [1:0] new_out12,
    output wire [1:0] new_out13,
    output wire [1:0] new_out14,
    output wire [1:0] new_out2,
    output wire [1:0] new_out3,
    output wire [1:0] new_out4,
    output wire [1:0] new_out7,
    output wire [2:0] new_out10,
    output wire [2:0] new_out11,
    output wire [2:0] new_out5,
    output wire [2:0] new_out6,
    output wire [2:0] new_out8,
    output wire [2:0] new_out9
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
wire w_060_;
wire w_061_;
wire w_062_;
wire w_063_;
wire w_064_;
wire w_065_;
wire w_066_;
wire w_067_;
wire w_068_;
wire w_069_;
wire w_070_;
wire w_071_;
wire w_072_;
wire w_073_;
wire w_074_;
wire w_075_;
wire w_076_;
wire w_077_;
wire w_078_;
wire w_079_;
wire w_080_;
wire w_081_;
wire w_082_;
wire w_083_;
wire w_084_;
wire w_085_;
wire w_086_;
wire w_087_;
wire w_088_;
wire w_089_;
wire w_090_;
wire w_091_;
wire w_092_;
wire w_093_;
wire w_094_;
wire w_095_;
wire w_096_;
wire w_097_;
wire w_098_;
wire w_099_;
wire w_100_;
wire w_101_;
wire w_102_;
wire w_103_;
wire w_104_;
wire w_105_;
wire w_106_;
wire w_107_;
wire w_108_;
wire w_109_;
wire w_110_;
wire w_111_;
wire w_112_;
wire w_113_;
wire w_114_;
wire w_115_;
wire w_116_;
wire w_117_;
wire w_118_;
wire w_119_;
wire w_120_;
wire w_121_;
wire w_122_;
wire w_123_;
wire w_124_;
wire w_125_;
wire w_126_;
wire w_127_;
wire w_128_;
wire w_129_;
wire w_130_;
wire w_131_;
wire w_132_;
wire w_133_;
wire w_134_;
wire w_135_;
wire w_136_;
wire w_137_;
wire w_138_;
wire w_139_;
wire w_140_;
wire w_141_;
wire w_142_;
wire w_143_;
wire w_144_;
wire w_145_;
wire w_146_;
wire w_147_;
wire w_148_;
wire w_149_;
wire w_150_;
wire w_151_;
wire w_152_;
wire w_153_;
wire w_154_;
wire w_155_;
wire w_156_;
wire w_157_;
wire w_158_;
wire w_159_;
wire w_160_;
wire w_161_;
wire w_162_;
wire w_163_;
wire w_164_;
wire w_165_;
wire w_166_;
wire w_167_;
wire w_168_;
wire w_169_;
wire w_170_;
wire w_171_;
wire w_172_;
wire w_173_;
wire w_174_;
wire w_175_;
wire w_176_;
wire w_177_;
wire w_178_;
wire w_179_;
wire w_180_;
wire w_181_;
wire w_182_;
wire w_183_;
wire w_184_;
wire w_185_;
wire w_186_;
wire w_187_;
wire w_188_;
wire w_189_;
wire w_190_;
wire w_191_;
wire w_192_;
wire w_193_;
wire w_194_;
wire w_195_;
wire w_196_;
wire w_197_;
wire w_198_;
wire w_199_;
wire w_200_;
wire w_201_;
wire w_202_;
wire w_203_;
wire w_204_;
wire w_205_;
wire w_206_;
wire w_207_;
wire w_208_;
wire w_209_;
wire w_210_;
wire w_211_;
wire w_212_;
wire w_213_;
wire w_214_;
wire w_215_;
wire w_216_;
wire w_217_;
wire w_218_;
wire w_219_;
wire w_220_;
wire w_221_;
wire w_222_;
wire w_223_;
wire w_224_;
wire w_225_;
wire w_226_;
wire w_227_;
wire w_228_;
wire w_229_;
wire w_230_;
wire w_231_;
wire w_232_;
wire w_233_;
wire w_234_;
wire w_235_;
wire w_236_;
wire w_237_;
wire w_238_;
wire w_239_;
wire w_240_;
wire w_241_;
wire w_242_;
wire w_243_;
wire w_244_;
wire w_245_;
wire w_246_;
wire w_247_;
wire w_248_;
wire w_249_;
wire w_250_;
wire w_251_;
wire w_252_;
wire w_253_;
wire w_254_;
wire w_255_;
wire w_256_;
wire w_257_;
wire w_258_;
wire w_259_;
wire w_260_;
wire w_261_;
wire w_262_;
wire w_263_;
wire w_264_;
wire w_265_;
wire w_266_;
wire w_267_;
wire w_268_;
wire w_269_;
wire w_270_;
wire w_271_;
wire w_272_;
wire w_273_;
wire w_274_;
wire w_275_;
wire w_276_;
wire w_277_;
wire w_278_;
wire w_279_;
wire w_280_;
wire w_281_;
wire w_282_;
wire w_283_;
wire w_284_;
wire w_285_;
wire w_286_;
wire w_287_;
wire w_288_;
wire w_289_;
wire w_290_;
wire w_291_;
wire w_292_;
wire w_293_;
wire w_294_;
wire w_295_;
wire w_296_;
wire w_297_;
wire w_298_;
wire w_299_;
wire w_300_;
wire w_301_;
wire w_302_;
wire w_303_;
wire w_304_;
wire w_305_;
wire w_306_;
wire w_307_;
wire w_308_;
wire w_309_;
wire w_310_;
wire w_311_;
wire w_312_;
wire w_313_;
wire w_314_;
wire w_315_;
wire w_316_;
wire w_317_;
wire w_318_;
wire w_319_;
wire w_320_;
wire w_321_;
wire w_322_;
wire w_323_;
wire w_324_;
wire w_325_;
wire w_326_;
wire w_327_;
wire w_328_;
wire w_329_;
wire w_330_;
wire w_331_;
wire w_332_;
wire w_333_;
wire w_334_;
wire w_335_;
wire w_336_;
wire w_337_;
wire w_338_;
wire w_339_;
wire w_340_;
wire w_341_;
wire w_342_;
wire w_343_;
wire w_344_;
wire w_345_;
wire w_346_;
wire w_347_;
wire w_348_;
wire w_349_;
wire w_350_;
wire w_351_;
wire w_352_;
wire w_353_;
wire w_354_;
nand (w_228_, new_in5[3], new_in4[3]);
nand (w_060_, w_216_, w_191_);
nand (w_154_, w_305_, w_194_);
xor (w_339_, new_in15[5], w_136_);
nand (w_343_, w_341_, w_169_);
nor (new_out8[0], w_233_, w_043_);
xor (w_169_, new_in10[5], w_092_);
not (w_159_, w_292_);
xor (w_269_, w_328_, w_311_);
and (w_021_, w_324_, w_002_);
not (w_247_, w_180_);
nand (w_132_, w_113_, w_293_);
nand (w_290_, new_in6[1], w_007_);
and (w_067_, new_in11[0], new_in2[0]);
nand (w_265_, w_010_, w_098_);
and (new_out2[1], w_292_, w_306_);
xor (w_283_, new_in14[6], new_in13[6]);
and (w_252_, w_254_, w_009_);
nand (w_212_, new_in15[3], w_218_);
nand (w_341_, w_168_, w_342_);
or (w_160_, w_306_, w_172_);
xor (w_007_, w_344_, w_337_);
nand (w_025_, w_266_, w_354_);
nand (w_106_, w_297_, w_241_);
xor (w_116_, new_in1[4], new_in12[4]);
xor (w_218_, w_310_, w_207_);
nand (w_034_, w_095_, w_025_);
nand (w_180_, w_350_, w_015_);
nand (w_249_, w_170_, w_022_);
xor (w_125_, w_346_, w_127_);
xor (w_262_, w_284_, w_032_);
nand (w_096_, new_in2[3], new_in11[3]);
xor (new_out4[0], w_269_, w_262_);
not (w_242_, w_091_);
xor (w_057_, new_in15[3], w_218_);
xor (w_030_, new_in10[4], w_089_);
xor (new_out3[1], w_179_, w_289_);
and (w_148_, new_in9[0], w_210_);
xor (w_042_, w_049_, w_234_);
xor (w_104_, new_in15[1], w_280_);
nand (w_209_, w_026_, w_352_);
not (w_293_, w_037_);
xor (w_182_, w_300_, w_213_);
xor (w_139_, new_in6[1], w_007_);
nand (w_317_, w_348_, w_215_);
nand (w_038_, w_250_, w_190_);
nand (w_020_, new_in10[5], w_092_);
nand (w_056_, w_310_, w_207_);
not (w_000_, w_016_);
nand (w_075_, new_in3[2], new_in8[2]);
xor (w_138_, w_148_, w_255_);
xor (w_257_, w_091_, w_162_);
xor (new_out13[1], w_307_, w_279_);
nand (w_121_, w_196_, w_330_);
xor (w_171_, new_in6[2], w_029_);
not (w_322_, w_019_);
xor (w_080_, w_268_, w_200_);
xor (w_179_, w_338_, w_079_);
nand (w_294_, w_265_, w_173_);
xor (w_137_, w_134_, w_339_);
xor (w_136_, w_340_, w_240_);
nand (w_033_, w_023_, w_245_);
not (w_331_, w_230_);
xor (w_246_, new_in10[1], w_059_);
xor (w_105_, new_in11[1], new_in2[1]);
xor (new_out9[2], w_313_, w_256_);
nand (w_022_, w_340_, w_240_);
xor (new_out1[0], new_in9[0], w_210_);
or (w_309_, w_176_, w_151_);
xor (w_264_, w_217_, w_076_);
nand (w_235_, new_in9[2], w_296_);
xor (w_352_, w_277_, w_257_);
xor (w_124_, w_321_, w_167_);
nand (w_185_, new_in9[3], w_014_);
nand (w_302_, w_321_, w_167_);
nand (w_338_, w_115_, w_329_);
nand (w_064_, w_348_, w_144_);
xor (w_337_, new_in8[1], new_in3[1]);
xor (w_200_, w_335_, w_267_);
or (w_351_, w_016_, w_179_);
xor (w_275_, new_in3[0], new_in8[0]);
nand (w_065_, w_117_, w_165_);
not (w_261_, new_out2[0]);
xor (w_276_, w_147_, w_111_);
xor (w_259_, w_150_, w_055_);
nand (w_354_, w_148_, w_255_);
nand (w_254_, new_in10[3], w_003_);
xor (w_190_, new_in13[1], new_in14[1]);
nand (w_054_, w_046_, w_267_);
nand (w_217_, w_183_, w_123_);
xor (w_127_, new_in5[3], new_in4[3]);
or (w_028_, w_201_, w_273_);
xor (w_213_, new_in5[2], new_in4[2]);
nand (w_073_, w_048_, w_027_);
and (w_243_, w_220_, w_072_);
nand (w_004_, w_075_, w_087_);
xor (w_188_, w_021_, w_074_);
xor (w_292_, w_110_, w_104_);
nand (w_141_, new_in15[1], w_280_);
xor (w_177_, w_157_, w_066_);
nand (w_345_, w_137_, w_093_);
nand (w_336_, w_081_, w_231_);
nand (w_014_, w_235_, w_034_);
nand (w_214_, w_353_, w_057_);
nand (w_187_, w_150_, w_042_);
nand (w_256_, w_209_, w_226_);
nand (w_081_, new_in13[5], new_in14[5]);
nand (w_224_, w_187_, w_069_);
xor (w_173_, w_211_, w_054_);
nand (w_157_, w_096_, w_056_);
nand (w_231_, w_326_, w_244_);
nand (w_326_, w_035_, w_154_);
not (w_135_, w_017_);
nand (w_277_, w_351_, w_178_);
xor (new_out7[0], w_001_, w_039_);
nand (w_175_, new_in7[3], w_125_);
and (w_314_, w_184_, w_192_);
xor (w_094_, new_in4[1], new_in5[1]);
xor (new_out4[1], w_352_, w_286_);
xor (w_176_, w_113_, w_037_);
nand (w_012_, w_091_, w_162_);
xor (w_274_, new_in1[2], new_in12[2]);
xor (w_145_, new_in15[2], w_264_);
and (w_250_, new_in13[0], new_in14[0]);
xor (w_319_, w_265_, w_173_);
nand (w_102_, w_219_, w_108_);
nand (w_288_, new_in8[1], new_in3[1]);
nand (w_103_, w_175_, w_085_);
nand (w_300_, w_045_, w_164_);
xor (w_167_, new_in1[3], new_in12[3]);
xor (w_108_, new_in10[6], w_291_);
nand (w_263_, w_053_, w_205_);
or (w_316_, w_181_, w_243_);
and (new_out8[2], w_215_, w_072_);
and (w_251_, new_in10[0], w_271_);
xor (w_047_, w_150_, w_306_);
and (w_344_, new_in3[0], new_in8[0]);
or (w_184_, w_276_, w_159_);
nand (w_048_, w_208_, w_124_);
xor (w_016_, w_229_, w_145_);
nand (w_123_, w_067_, w_105_);
xor (w_072_, w_172_, w_086_);
nand (w_156_, new_in10[1], w_059_);
xor (w_074_, w_222_, w_253_);
nand (w_186_, new_in15[5], w_136_);
not (w_008_, w_297_);
not (w_301_, w_137_);
or (w_206_, w_301_, w_303_);
nand (w_036_, new_in5[2], new_in4[2]);
nand (w_324_, w_319_, w_114_);
nand (w_043_, w_034_, w_051_);
nand (w_312_, new_in7[1], w_083_);
not (w_287_, new_in6[0]);
and (w_197_, w_263_, w_140_);
xor (w_083_, w_199_, w_094_);
nand (w_321_, w_327_, w_248_);
xor (new_out13[0], new_out1[1], w_348_);
nand (w_340_, w_295_, w_133_);
and (w_061_, w_019_, w_155_);
xor (w_129_, w_068_, w_247_);
xor (w_349_, w_281_, w_032_);
xor (w_162_, w_353_, w_057_);
xor (w_194_, new_in14[4], new_in13[4]);
nand (w_011_, w_186_, w_166_);
or (w_146_, new_in9[4], w_204_);
xor (w_303_, w_219_, w_108_);
xor (w_181_, w_126_, w_013_);
xor (w_111_, new_in10[2], w_071_);
not (w_281_, new_out1[1]);
xor (new_out6[0], w_276_, w_000_);
or (w_193_, w_230_, w_239_);
xor (w_291_, w_336_, w_283_);
nand (w_023_, w_118_, w_065_);
xor (new_out10[0], w_345_, w_259_);
xor (new_out5[2], w_044_, w_047_);
nand (w_219_, w_020_, w_343_);
xor (w_112_, w_026_, w_352_);
xor (w_273_, w_129_, w_215_);
xor (w_245_, new_in13[3], new_in14[3]);
xor (w_126_, w_319_, w_114_);
nand (w_329_, w_147_, w_111_);
nand (w_031_, w_217_, w_076_);
nand (w_226_, w_121_, w_112_);
xor (w_306_, w_261_, w_237_);
and (new_out2[0], w_068_, w_180_);
and (w_203_, w_282_, w_316_);
nand (w_198_, w_129_, w_349_);
xor (w_109_, w_090_, w_320_);
and (w_107_, new_in6[0], w_275_);
nand (w_260_, new_in6[2], w_029_);
nand (w_236_, w_298_, w_302_);
nand (w_327_, new_in1[2], new_in12[2]);
nand (w_045_, new_in4[1], new_in5[1]);
nand (w_024_, w_049_, w_234_);
xor (w_268_, w_249_, w_011_);
xor (w_091_, w_252_, w_030_);
nand (w_098_, w_278_, w_080_);
xor (new_out10[1], w_061_, w_334_);
xor (w_086_, w_176_, w_151_);
and (w_332_, w_196_, w_227_);
nand (w_168_, new_in10[4], w_089_);
xor (w_286_, w_325_, w_320_);
nand (w_267_, w_299_, w_102_);
xor (w_325_, w_149_, w_171_);
or (w_015_, w_251_, w_246_);
nand (w_118_, new_in14[2], new_in13[2]);
xor (w_220_, w_058_, w_253_);
and (w_114_, w_224_, w_253_);
nand (w_149_, w_290_, w_006_);
nand (w_069_, w_174_, w_258_);
xor (w_032_, w_107_, w_139_);
nand (w_046_, w_163_, w_153_);
nand (w_350_, w_251_, w_246_);
xor (w_232_, w_287_, w_275_);
and (w_297_, new_in7[0], w_062_);
nand (w_134_, w_223_, w_063_);
xor (w_241_, new_in7[1], w_083_);
nand (w_050_, w_141_, w_189_);
xor (w_237_, w_276_, w_159_);
nand (w_009_, w_338_, w_079_);
xor (w_271_, new_in13[0], new_in14[0]);
xor (new_out3[0], w_276_, w_233_);
nand (w_315_, w_288_, w_005_);
xor (w_013_, w_109_, w_042_);
nand (w_006_, w_107_, w_139_);
nand (w_005_, w_344_, w_337_);
nand (w_238_, w_313_, w_256_);
nand (w_227_, w_269_, w_109_);
xor (w_313_, w_215_, w_086_);
xor (new_out11[2], w_188_, w_203_);
nand (w_087_, w_315_, w_308_);
nand (w_128_, w_228_, w_225_);
and (w_334_, w_197_, w_268_);
nand (w_270_, w_215_, w_086_);
nand (w_130_, w_052_, w_101_);
and (w_307_, new_out1[1], w_348_);
and (w_211_, w_249_, w_011_);
xor (w_099_, w_082_, w_078_);
nand (w_330_, w_122_, w_227_);
nand (new_out12[1], w_180_, w_109_);
nand (w_084_, new_in15[2], w_264_);
nand (w_122_, w_160_, w_143_);
xor (new_out14[1], w_272_, w_138_);
xor (w_207_, new_in2[3], new_in11[3]);
nand (w_035_, new_in14[4], new_in13[4]);
not (w_026_, w_222_);
xor (new_out5[1], w_201_, w_273_);
xor (w_284_, w_008_, w_241_);
nand (w_147_, w_156_, w_350_);
xor (w_003_, w_023_, w_245_);
xor (w_289_, w_144_, w_352_);
nand (w_311_, w_184_, w_192_);
xor (w_272_, w_122_, w_332_);
and (w_199_, new_in4[0], new_in5[0]);
xor (w_308_, new_in3[2], new_in8[2]);
nand (w_305_, w_347_, w_033_);
not (w_040_, w_220_);
or (w_208_, new_in9[3], w_014_);
nand (w_101_, w_285_, w_088_);
nand (w_278_, w_206_, w_024_);
xor (w_092_, w_326_, w_244_);
not (w_333_, w_013_);
nand (w_077_, w_300_, w_213_);
nand (w_163_, new_in14[6], new_in13[6]);
xor (w_066_, new_in2[4], new_in11[4]);
xor (w_240_, new_in11[5], new_in2[5]);
nand (w_295_, new_in2[4], new_in11[4]);
nand (w_155_, w_150_, w_055_);
xor (new_out7[1], new_out9[2], w_318_);
nand (w_153_, w_336_, w_283_);
or (w_196_, w_269_, w_109_);
nand (w_049_, w_132_, w_309_);
nand (w_225_, w_346_, w_127_);
xor (new_out9[1], w_322_, w_001_);
xor (w_082_, w_306_, w_172_);
xor (w_029_, w_315_, w_308_);
xor (w_100_, new_in7[3], w_125_);
nor (new_out8[1], w_135_, w_289_);
nand (w_183_, new_in11[1], new_in2[1]);
nand (w_310_, w_202_, w_031_);
nand (w_133_, w_157_, w_066_);
nand (w_119_, w_277_, w_257_);
xor (w_165_, new_in14[2], new_in13[2]);
xor (w_071_, w_117_, w_165_);
nand (w_158_, w_260_, w_142_);
xor (new_out5[0], w_230_, w_222_);
nand (w_192_, new_out2[0], w_237_);
xor (w_230_, new_in10[0], w_271_);
nand (w_189_, w_110_, w_104_);
and (w_002_, w_131_, w_294_);
nand (w_019_, w_004_, w_158_);
not (w_229_, w_050_);
xor (w_055_, w_004_, w_158_);
nand (w_248_, w_161_, w_274_);
nand (new_out12[0], w_331_, w_172_);
xor (w_172_, w_284_, w_325_);
xor (w_210_, new_in1[0], new_in12[0]);
xor (w_088_, new_in7[2], w_182_);
or (w_178_, w_328_, w_314_);
not (w_335_, w_046_);
and (w_039_, w_292_, w_138_);
nand (w_304_, w_050_, w_145_);
and (w_078_, w_198_, w_097_);
nand (w_142_, w_149_, w_171_);
xor (w_348_, w_068_, w_180_);
nand (w_342_, w_323_, w_030_);
nand (w_115_, new_in10[2], w_071_);
xor (new_out6[1], w_179_, w_162_);
nand (w_299_, new_in10[6], w_291_);
nand (w_298_, new_in1[3], new_in12[3]);
nand (w_353_, w_084_, w_304_);
nand (w_097_, w_064_, w_193_);
and (w_151_, w_012_, w_119_);
xor (new_out9[0], w_055_, w_272_);
not (w_144_, w_349_);
xor (w_113_, w_120_, w_018_);
xor (w_079_, new_in10[3], w_003_);
xor (w_244_, new_in13[5], new_in14[5]);
xor (w_279_, w_306_, w_284_);
nand (w_053_, new_in1[4], new_in12[4]);
nand (w_285_, w_312_, w_106_);
xor (w_070_, new_in11[0], new_in2[0]);
nand (w_170_, new_in11[5], new_in2[5]);
xor (w_239_, new_out1[0], w_232_);
and (w_150_, w_128_, w_103_);
and (w_044_, w_317_, w_028_);
or (w_051_, w_095_, w_025_);
xor (w_280_, w_067_, w_105_);
nand (w_346_, w_036_, w_077_);
xor (w_018_, new_in15[4], w_177_);
nand (w_085_, w_130_, w_100_);
xor (w_089_, w_305_, w_194_);
or (w_201_, w_230_, w_222_);
and (w_216_, new_in1[0], new_in12[0]);
xor (w_320_, w_285_, w_088_);
xor (w_215_, w_128_, w_103_);
nor (w_318_, w_016_, w_043_);
xor (w_037_, w_341_, w_169_);
xor (w_222_, w_019_, w_017_);
nand (w_117_, w_195_, w_038_);
nand (w_266_, new_in9[1], w_041_);
xor (w_233_, w_239_, w_269_);
nand (w_202_, new_in2[2], new_in11[2]);
xor (w_296_, w_161_, w_274_);
xor (w_234_, w_301_, w_303_);
xor (w_204_, w_236_, w_116_);
xor (new_out14[0], new_out1[0], w_099_);
xor (w_017_, w_130_, w_100_);
nand (w_143_, w_082_, w_078_);
xor (w_255_, new_in9[1], w_041_);
xor (new_out11[0], w_040_, w_072_);
xor (new_out11[1], w_181_, w_243_);
nand (w_161_, w_221_, w_060_);
xor (w_191_, new_in12[1], new_in1[1]);
and (w_140_, w_146_, w_073_);
nand (w_282_, w_126_, w_333_);
nand (w_195_, new_in13[1], new_in14[1]);
xor (w_328_, w_000_, w_179_);
xor (w_059_, w_250_, w_190_);
nand (w_166_, w_134_, w_339_);
xor (new_out6[2], w_242_, w_113_);
nand (w_258_, w_270_, w_238_);
xor (w_093_, w_263_, w_140_);
nand (w_205_, w_236_, w_116_);
xor (w_001_, w_121_, w_112_);
and (w_027_, w_152_, w_185_);
nand (w_120_, w_212_, w_214_);
xor (w_068_, new_in15[0], w_070_);
nand (w_063_, w_120_, w_018_);
nand (w_052_, new_in7[2], w_182_);
nand (w_323_, w_254_, w_009_);
xor (w_041_, w_216_, w_191_);
xor (new_out1[1], new_in7[0], w_062_);
or (w_174_, w_150_, w_042_);
xor (w_095_, new_in9[2], w_296_);
nand (w_164_, w_199_, w_094_);
nand (w_223_, new_in15[4], w_177_);
xor (w_253_, w_278_, w_080_);
xor (w_076_, new_in2[2], new_in11[2]);
xor (w_062_, new_in4[0], new_in5[0]);
nand (w_131_, w_211_, w_054_);
not (w_090_, w_055_);
nand (w_347_, new_in13[3], new_in14[3]);
nand (w_152_, new_in9[4], w_204_);
and (w_110_, new_in15[0], w_070_);
nand (w_010_, w_268_, w_200_);
nand (w_221_, new_in12[1], new_in1[1]);
not (w_058_, w_224_);
buf (new_out10[2], 1'h1);
endmodule
