module sub_module1(
    input wire in1,
    input wire in2,
    input wire in3,
    input wire in4,
    input wire in5,
    input wire in6,
    input wire in7,
    input wire in8,
    input wire in9,
    input wire in10,
    input wire in11,
    input wire in12,
    input wire in13,
    input wire in14,
    input wire in15,
    input wire in16,
    output wire out1,
    output wire out2,
    output wire out3,
    output wire out4,
    output wire out5,
    output wire out6,
    output wire out7,
    output wire out8,
    output wire out9,
    output wire out10
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
wire w_060_;
wire w_061_;
wire w_062_;
wire w_063_;
wire w_064_;
wire w_065_;
wire w_066_;
wire w_067_;
wire w_068_;
wire w_069_;
wire w_070_;
wire w_071_;
wire w_072_;
wire w_073_;
wire w_074_;
wire w_075_;
wire w_076_;
wire w_077_;
wire w_078_;
wire w_079_;
wire w_080_;
wire w_081_;
wire w_082_;
wire w_083_;
wire w_084_;
wire w_085_;
wire w_086_;
wire w_087_;
wire w_088_;
wire w_089_;
wire w_090_;
wire w_091_;
wire w_092_;
wire w_093_;
wire w_094_;
wire w_095_;
wire w_096_;
wire w_097_;
wire w_098_;
wire w_099_;
wire w_100_;
wire w_101_;
wire w_102_;
wire w_103_;
wire w_104_;
wire w_105_;
wire w_106_;
wire w_107_;
or (w_036_, w_044_, w_076_);
not (w_092_, w_062_);
or (w_096_, w_029_, w_083_);
not (w_025_, in2);
not (w_107_, in1);
not (w_070_, w_022_);
not (w_021_, w_088_);
or (w_023_, in4, in8);
and (w_007_, w_045_, w_026_);
or (w_027_, w_067_, w_007_);
and (out10, w_104_, w_057_);
or (w_078_, w_045_, w_026_);
or (w_002_, in12, in6);
and (w_067_, w_071_, w_074_);
or (w_034_, w_000_, w_087_);
or (w_006_, in8, w_028_);
and (w_068_, in1, in9);
or (w_104_, w_040_, w_103_);
or (w_062_, w_093_, w_051_);
not (out1, w_099_);
not (w_105_, w_058_);
or (w_057_, w_096_, w_060_);
and (w_058_, in15, in16);
or (out2, w_055_, w_086_);
or (w_094_, w_006_, w_056_);
not (w_085_, w_036_);
or (w_074_, in3, in4);
and (w_040_, w_054_, w_016_);
not (w_049_, in12);
and (w_030_, w_034_, w_096_);
and (w_048_, w_099_, w_046_);
and (out9, w_019_, w_096_);
or (w_063_, in12, w_053_);
or (w_099_, w_037_, w_032_);
and (w_084_, in3, in11);
or (w_009_, in10, in2);
or (w_031_, in6, w_004_);
and (w_052_, in6, w_004_);
not (w_015_, w_061_);
or (w_080_, w_065_, w_003_);
and (w_079_, w_027_, w_093_);
not (w_005_, out4);
or (w_060_, w_038_, w_048_);
and (w_056_, w_106_, w_079_);
and (w_032_, w_006_, w_027_);
not (w_024_, in8);
and (out7, w_090_, w_094_);
or (w_097_, w_070_, w_058_);
and (w_086_, w_006_, w_020_);
and (w_095_, w_106_, w_093_);
or (w_076_, w_009_, w_072_);
and (w_017_, in13, in15);
not (out3, w_046_);
and (w_045_, in1, w_025_);
or (w_046_, w_095_, w_021_);
and (w_012_, w_005_, w_062_);
and (w_039_, w_024_, w_050_);
and (w_001_, w_039_, out4);
and (w_053_, w_102_, w_010_);
and (w_018_, w_091_, w_073_);
or (w_082_, w_071_, w_074_);
and (w_010_, in9, in10);
not (w_064_, w_052_);
and (w_103_, w_011_, w_100_);
and (w_091_, w_084_, w_017_);
and (w_073_, w_004_, w_068_);
and (w_061_, in13, in14);
not (w_013_, w_018_);
not (w_090_, w_019_);
or (w_050_, w_101_, w_052_);
not (w_059_, w_033_);
and (w_106_, w_098_, w_097_);
and (w_019_, w_006_, w_056_);
not (w_102_, in11);
or (w_098_, w_081_, w_061_);
or (out6, w_001_, w_042_);
and (w_014_, w_096_, w_089_);
and (w_043_, out4, w_092_);
not (w_003_, in10);
or (out8, w_043_, w_012_);
and (w_083_, w_018_, w_085_);
or (w_022_, in15, in16);
or (w_051_, w_006_, w_027_);
or (w_072_, in14, in16);
and (w_069_, w_035_, w_020_);
or (w_044_, w_023_, w_002_);
or (w_066_, in13, in14);
or (out4, w_030_, w_075_);
not (w_065_, in9);
and (w_087_, w_022_, w_105_);
not (w_026_, w_074_);
or (w_071_, w_107_, in2);
and (w_004_, in5, in7);
not (w_101_, w_031_);
or (w_047_, in11, w_080_);
or (w_016_, w_013_, w_036_);
or (w_089_, w_079_, w_069_);
and (w_028_, w_031_, w_064_);
or (w_093_, w_041_, w_063_);
or (w_008_, w_102_, w_010_);
and (w_035_, w_078_, w_082_);
and (w_041_, in11, w_080_);
and (w_042_, w_006_, w_005_);
and (w_077_, w_049_, w_008_);
and (w_037_, w_039_, w_035_);
or (w_054_, w_018_, w_085_);
or (w_088_, w_106_, w_093_);
or (w_100_, out1, out3);
and (w_000_, w_066_, w_015_);
and (w_038_, out1, out3);
and (w_029_, w_013_, w_036_);
and (w_055_, w_039_, w_093_);
or (w_033_, w_096_, w_089_);
not (w_081_, w_066_);
or (out5, w_014_, w_059_);
or (w_011_, w_099_, w_046_);
and (w_020_, w_047_, w_077_);
and (w_075_, w_106_, w_040_);
endmodule

module sub_module2(
    input wire [5:0] in1,
    input wire [5:0] in2,
    input wire [5:0] in3,
    input wire [5:0] in4,
    input wire [5:0] in5,
    input wire [5:0] in6,
    input wire [5:0] in7,
    input wire [5:0] in8,
    input wire [7:0] in9,
    input wire [7:0] in10,
    input wire [7:0] in11,
    input wire [7:0] in12,
    input wire [7:0] in13,
    input wire [7:0] in14,
    input wire [7:0] in15,
    input wire [7:0] in16,
    output wire [5:0] out1,
    output wire [5:0] out2,
    output wire [5:0] out3,
    output wire [5:0] out4,
    output wire [5:0] out5,
    output wire [5:0] out6,
    output wire [5:0] out7,
    output wire [5:0] out8,
    output wire [5:0] out9,
    output wire [5:0] out10,
    output wire [5:0] out11,
    output wire [5:0] out12,
    output wire [7:0] out13,
    output wire [7:0] out14,
    output wire [7:0] out15,
    output wire [7:0] out16,
    output wire [7:0] out17,
    output wire [7:0] out18,
    output wire [7:0] out19,
    output wire [7:0] out20,
    output wire [7:0] out21,
    output wire [7:0] out22,
    output wire [7:0] out23,
    output wire [7:0] out24
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
wire w_0945_;
wire w_0946_;
wire w_0947_;
wire w_0948_;
wire w_0949_;
wire w_0950_;
wire w_0951_;
wire w_0952_;
wire w_0953_;
wire w_0954_;
wire w_0955_;
wire w_0956_;
wire w_0957_;
wire w_0958_;
wire w_0959_;
wire w_0960_;
wire w_0961_;
wire w_0962_;
wire w_0963_;
wire w_0964_;
wire w_0965_;
wire w_0966_;
wire w_0967_;
wire w_0968_;
wire w_0969_;
wire w_0970_;
wire w_0971_;
wire w_0972_;
wire w_0973_;
wire w_0974_;
wire w_0975_;
wire w_0976_;
wire w_0977_;
wire w_0978_;
wire w_0979_;
wire w_0980_;
wire w_0981_;
wire w_0982_;
wire w_0983_;
wire w_0984_;
wire w_0985_;
wire w_0986_;
wire w_0987_;
wire w_0988_;
wire w_0989_;
wire w_0990_;
wire w_0991_;
wire w_0992_;
wire w_0993_;
wire w_0994_;
wire w_0995_;
wire w_0996_;
wire w_0997_;
wire w_0998_;
wire w_0999_;
wire w_1000_;
wire w_1001_;
wire w_1002_;
wire w_1003_;
wire w_1004_;
wire w_1005_;
wire w_1006_;
wire w_1007_;
wire w_1008_;
wire w_1009_;
wire w_1010_;
wire w_1011_;
wire w_1012_;
wire w_1013_;
wire w_1014_;
wire w_1015_;
wire w_1016_;
wire w_1017_;
wire w_1018_;
wire w_1019_;
wire w_1020_;
wire w_1021_;
wire w_1022_;
wire w_1023_;
wire w_1024_;
wire w_1025_;
wire w_1026_;
wire w_1027_;
wire w_1028_;
wire w_1029_;
wire w_1030_;
wire w_1031_;
wire w_1032_;
wire w_1033_;
wire w_1034_;
wire w_1035_;
wire w_1036_;
wire w_1037_;
wire w_1038_;
wire w_1039_;
wire w_1040_;
wire w_1041_;
wire w_1042_;
wire w_1043_;
wire w_1044_;
wire w_1045_;
wire w_1046_;
wire w_1047_;
wire w_1048_;
wire w_1049_;
wire w_1050_;
wire w_1051_;
wire w_1052_;
wire w_1053_;
wire w_1054_;
wire w_1055_;
wire w_1056_;
wire w_1057_;
wire w_1058_;
wire w_1059_;
wire w_1060_;
wire w_1061_;
wire w_1062_;
wire w_1063_;
wire w_1064_;
wire w_1065_;
wire w_1066_;
wire w_1067_;
wire w_1068_;
wire w_1069_;
wire w_1070_;
wire w_1071_;
wire w_1072_;
wire w_1073_;
wire w_1074_;
wire w_1075_;
wire w_1076_;
wire w_1077_;
wire w_1078_;
wire w_1079_;
wire w_1080_;
wire w_1081_;
wire w_1082_;
wire w_1083_;
wire w_1084_;
wire w_1085_;
wire w_1086_;
wire w_1087_;
wire w_1088_;
wire w_1089_;
wire w_1090_;
wire w_1091_;
wire w_1092_;
wire w_1093_;
wire w_1094_;
wire w_1095_;
wire w_1096_;
wire w_1097_;
wire w_1098_;
wire w_1099_;
wire w_1100_;
wire w_1101_;
wire w_1102_;
wire w_1103_;
wire w_1104_;
wire w_1105_;
wire w_1106_;
wire w_1107_;
wire w_1108_;
wire w_1109_;
wire w_1110_;
wire w_1111_;
wire w_1112_;
wire w_1113_;
wire w_1114_;
wire w_1115_;
wire w_1116_;
wire w_1117_;
wire w_1118_;
wire w_1119_;
wire w_1120_;
wire w_1121_;
wire w_1122_;
wire w_1123_;
wire w_1124_;
wire w_1125_;
wire w_1126_;
wire w_1127_;
wire w_1128_;
wire w_1129_;
wire w_1130_;
wire w_1131_;
wire w_1132_;
wire w_1133_;
wire w_1134_;
wire w_1135_;
wire w_1136_;
wire w_1137_;
wire w_1138_;
wire w_1139_;
wire w_1140_;
wire w_1141_;
wire w_1142_;
wire w_1143_;
wire w_1144_;
wire w_1145_;
wire w_1146_;
wire w_1147_;
wire w_1148_;
wire w_1149_;
wire w_1150_;
wire w_1151_;
wire w_1152_;
wire w_1153_;
wire w_1154_;
wire w_1155_;
wire w_1156_;
wire w_1157_;
wire w_1158_;
wire w_1159_;
wire w_1160_;
wire w_1161_;
wire w_1162_;
wire w_1163_;
wire w_1164_;
wire w_1165_;
wire w_1166_;
wire w_1167_;
wire w_1168_;
wire w_1169_;
wire w_1170_;
wire w_1171_;
wire w_1172_;
wire w_1173_;
wire w_1174_;
wire w_1175_;
wire w_1176_;
wire w_1177_;
wire w_1178_;
wire w_1179_;
wire w_1180_;
wire w_1181_;
wire w_1182_;
wire w_1183_;
wire w_1184_;
wire w_1185_;
wire w_1186_;
wire w_1187_;
wire w_1188_;
wire w_1189_;
wire w_1190_;
wire w_1191_;
wire w_1192_;
wire w_1193_;
wire w_1194_;
wire w_1195_;
wire w_1196_;
wire w_1197_;
wire w_1198_;
wire w_1199_;
wire w_1200_;
wire w_1201_;
wire w_1202_;
wire w_1203_;
wire w_1204_;
wire w_1205_;
wire w_1206_;
wire w_1207_;
wire w_1208_;
wire w_1209_;
wire w_1210_;
wire w_1211_;
wire w_1212_;
wire w_1213_;
wire w_1214_;
wire w_1215_;
wire w_1216_;
wire w_1217_;
wire w_1218_;
wire w_1219_;
wire w_1220_;
wire w_1221_;
wire w_1222_;
wire w_1223_;
wire w_1224_;
wire w_1225_;
wire w_1226_;
wire w_1227_;
wire w_1228_;
wire w_1229_;
wire w_1230_;
wire w_1231_;
wire w_1232_;
wire w_1233_;
wire w_1234_;
wire w_1235_;
wire w_1236_;
wire w_1237_;
wire w_1238_;
wire w_1239_;
wire w_1240_;
wire w_1241_;
wire w_1242_;
wire w_1243_;
wire w_1244_;
wire w_1245_;
wire w_1246_;
wire w_1247_;
wire w_1248_;
wire w_1249_;
wire w_1250_;
wire w_1251_;
wire w_1252_;
wire w_1253_;
wire w_1254_;
wire w_1255_;
wire w_1256_;
wire w_1257_;
wire w_1258_;
wire w_1259_;
wire w_1260_;
wire w_1261_;
wire w_1262_;
wire w_1263_;
wire w_1264_;
wire w_1265_;
wire w_1266_;
wire w_1267_;
wire w_1268_;
wire w_1269_;
wire w_1270_;
wire w_1271_;
wire w_1272_;
wire w_1273_;
wire w_1274_;
wire w_1275_;
wire w_1276_;
wire w_1277_;
wire w_1278_;
wire w_1279_;
wire w_1280_;
wire w_1281_;
wire w_1282_;
wire w_1283_;
wire w_1284_;
wire w_1285_;
wire w_1286_;
wire w_1287_;
wire w_1288_;
wire w_1289_;
wire w_1290_;
wire w_1291_;
wire w_1292_;
wire w_1293_;
wire w_1294_;
wire w_1295_;
wire w_1296_;
wire w_1297_;
wire w_1298_;
wire w_1299_;
wire w_1300_;
wire w_1301_;
wire w_1302_;
wire w_1303_;
wire w_1304_;
wire w_1305_;
wire w_1306_;
wire w_1307_;
wire w_1308_;
wire w_1309_;
wire w_1310_;
wire w_1311_;
wire w_1312_;
wire w_1313_;
wire w_1314_;
wire w_1315_;
wire w_1316_;
wire w_1317_;
wire w_1318_;
wire w_1319_;
wire w_1320_;
wire w_1321_;
wire w_1322_;
wire w_1323_;
wire w_1324_;
wire w_1325_;
wire w_1326_;
wire w_1327_;
wire w_1328_;
wire w_1329_;
wire w_1330_;
wire w_1331_;
wire w_1332_;
wire w_1333_;
wire w_1334_;
wire w_1335_;
wire w_1336_;
wire w_1337_;
wire w_1338_;
wire w_1339_;
wire w_1340_;
wire w_1341_;
wire w_1342_;
wire w_1343_;
wire w_1344_;
wire w_1345_;
wire w_1346_;
wire w_1347_;
wire w_1348_;
wire w_1349_;
wire w_1350_;
wire w_1351_;
wire w_1352_;
wire w_1353_;
wire w_1354_;
wire w_1355_;
wire w_1356_;
wire w_1357_;
wire w_1358_;
wire w_1359_;
wire w_1360_;
wire w_1361_;
wire w_1362_;
wire w_1363_;
wire w_1364_;
wire w_1365_;
wire w_1366_;
wire w_1367_;
wire w_1368_;
wire w_1369_;
wire w_1370_;
wire w_1371_;
wire w_1372_;
wire w_1373_;
wire w_1374_;
wire w_1375_;
wire w_1376_;
wire w_1377_;
wire w_1378_;
wire w_1379_;
wire w_1380_;
wire w_1381_;
wire w_1382_;
wire w_1383_;
wire w_1384_;
wire w_1385_;
wire w_1386_;
wire w_1387_;
wire w_1388_;
wire w_1389_;
wire w_1390_;
wire w_1391_;
wire w_1392_;
wire w_1393_;
wire w_1394_;
wire w_1395_;
wire w_1396_;
wire w_1397_;
wire w_1398_;
wire w_1399_;
wire w_1400_;
wire w_1401_;
wire w_1402_;
wire w_1403_;
wire w_1404_;
wire w_1405_;
wire w_1406_;
wire w_1407_;
wire w_1408_;
wire w_1409_;
wire w_1410_;
wire w_1411_;
wire w_1412_;
wire w_1413_;
wire w_1414_;
wire w_1415_;
wire w_1416_;
wire w_1417_;
wire w_1418_;
wire w_1419_;
wire w_1420_;
wire w_1421_;
wire w_1422_;
wire w_1423_;
wire w_1424_;
wire w_1425_;
wire w_1426_;
wire w_1427_;
wire w_1428_;
wire w_1429_;
wire w_1430_;
wire w_1431_;
wire w_1432_;
wire w_1433_;
wire w_1434_;
wire w_1435_;
wire w_1436_;
wire w_1437_;
wire w_1438_;
wire w_1439_;
wire w_1440_;
wire w_1441_;
wire w_1442_;
wire w_1443_;
wire w_1444_;
wire w_1445_;
wire w_1446_;
wire w_1447_;
wire w_1448_;
wire w_1449_;
wire w_1450_;
wire w_1451_;
wire w_1452_;
wire w_1453_;
wire w_1454_;
wire w_1455_;
wire w_1456_;
wire w_1457_;
wire w_1458_;
wire w_1459_;
wire w_1460_;
wire w_1461_;
wire w_1462_;
wire w_1463_;
wire w_1464_;
wire w_1465_;
wire w_1466_;
wire w_1467_;
wire w_1468_;
wire w_1469_;
wire w_1470_;
wire w_1471_;
wire w_1472_;
wire w_1473_;
wire w_1474_;
wire w_1475_;
wire w_1476_;
wire w_1477_;
wire w_1478_;
wire w_1479_;
wire w_1480_;
wire w_1481_;
wire w_1482_;
wire w_1483_;
wire w_1484_;
wire w_1485_;
wire w_1486_;
wire w_1487_;
wire w_1488_;
wire w_1489_;
wire w_1490_;
wire w_1491_;
wire w_1492_;
wire w_1493_;
wire w_1494_;
wire w_1495_;
wire w_1496_;
wire w_1497_;
wire w_1498_;
wire w_1499_;
wire w_1500_;
wire w_1501_;
wire w_1502_;
wire w_1503_;
wire w_1504_;
wire w_1505_;
wire w_1506_;
wire w_1507_;
wire w_1508_;
wire w_1509_;
wire w_1510_;
wire w_1511_;
wire w_1512_;
wire w_1513_;
wire w_1514_;
wire w_1515_;
wire w_1516_;
wire w_1517_;
wire w_1518_;
wire w_1519_;
wire w_1520_;
wire w_1521_;
wire w_1522_;
wire w_1523_;
wire w_1524_;
wire w_1525_;
wire w_1526_;
wire w_1527_;
wire w_1528_;
wire w_1529_;
wire w_1530_;
wire w_1531_;
wire w_1532_;
wire w_1533_;
wire w_1534_;
wire w_1535_;
wire w_1536_;
wire w_1537_;
wire w_1538_;
wire w_1539_;
wire w_1540_;
wire w_1541_;
wire w_1542_;
wire w_1543_;
wire w_1544_;
wire w_1545_;
wire w_1546_;
wire w_1547_;
wire w_1548_;
wire w_1549_;
wire w_1550_;
wire w_1551_;
wire w_1552_;
wire w_1553_;
wire w_1554_;
wire w_1555_;
wire w_1556_;
wire w_1557_;
wire w_1558_;
wire w_1559_;
wire w_1560_;
wire w_1561_;
wire w_1562_;
wire w_1563_;
wire w_1564_;
wire w_1565_;
wire w_1566_;
wire w_1567_;
wire w_1568_;
wire w_1569_;
wire w_1570_;
wire w_1571_;
wire w_1572_;
wire w_1573_;
wire w_1574_;
wire w_1575_;
wire w_1576_;
wire w_1577_;
wire w_1578_;
wire w_1579_;
wire w_1580_;
wire w_1581_;
wire w_1582_;
wire w_1583_;
wire w_1584_;
wire w_1585_;
wire w_1586_;
wire w_1587_;
wire w_1588_;
wire w_1589_;
wire w_1590_;
wire w_1591_;
wire w_1592_;
wire w_1593_;
wire w_1594_;
wire w_1595_;
wire w_1596_;
wire w_1597_;
wire w_1598_;
wire w_1599_;
wire w_1600_;
wire w_1601_;
wire w_1602_;
wire w_1603_;
wire w_1604_;
wire w_1605_;
wire w_1606_;
wire w_1607_;
wire w_1608_;
wire w_1609_;
wire w_1610_;
wire w_1611_;
wire w_1612_;
wire w_1613_;
wire w_1614_;
wire w_1615_;
wire w_1616_;
wire w_1617_;
wire w_1618_;
wire w_1619_;
wire w_1620_;
wire w_1621_;
wire w_1622_;
wire w_1623_;
wire w_1624_;
wire w_1625_;
wire w_1626_;
wire w_1627_;
wire w_1628_;
wire w_1629_;
wire w_1630_;
wire w_1631_;
wire w_1632_;
wire w_1633_;
wire w_1634_;
wire w_1635_;
wire w_1636_;
wire w_1637_;
wire w_1638_;
wire w_1639_;
wire w_1640_;
wire w_1641_;
wire w_1642_;
wire w_1643_;
wire w_1644_;
wire w_1645_;
wire w_1646_;
wire w_1647_;
wire w_1648_;
wire w_1649_;
wire w_1650_;
wire w_1651_;
wire w_1652_;
wire w_1653_;
wire w_1654_;
wire w_1655_;
wire w_1656_;
wire w_1657_;
wire w_1658_;
wire w_1659_;
wire w_1660_;
wire w_1661_;
wire w_1662_;
wire w_1663_;
wire w_1664_;
wire w_1665_;
wire w_1666_;
wire w_1667_;
wire w_1668_;
wire w_1669_;
wire w_1670_;
wire w_1671_;
wire w_1672_;
wire w_1673_;
wire w_1674_;
wire w_1675_;
wire w_1676_;
wire w_1677_;
wire w_1678_;
wire w_1679_;
wire w_1680_;
wire w_1681_;
wire w_1682_;
wire w_1683_;
wire w_1684_;
wire w_1685_;
wire w_1686_;
wire w_1687_;
wire w_1688_;
wire w_1689_;
wire w_1690_;
wire w_1691_;
wire w_1692_;
wire w_1693_;
wire w_1694_;
wire w_1695_;
wire w_1696_;
wire w_1697_;
wire w_1698_;
wire w_1699_;
wire w_1700_;
wire w_1701_;
wire w_1702_;
wire w_1703_;
wire w_1704_;
wire w_1705_;
wire w_1706_;
wire w_1707_;
wire w_1708_;
wire w_1709_;
wire w_1710_;
wire w_1711_;
wire w_1712_;
wire w_1713_;
wire w_1714_;
wire w_1715_;
wire w_1716_;
wire w_1717_;
wire w_1718_;
wire w_1719_;
wire w_1720_;
wire w_1721_;
wire w_1722_;
wire w_1723_;
wire w_1724_;
wire w_1725_;
wire w_1726_;
wire w_1727_;
wire w_1728_;
wire w_1729_;
wire w_1730_;
wire w_1731_;
wire w_1732_;
wire w_1733_;
wire w_1734_;
wire w_1735_;
wire w_1736_;
wire w_1737_;
wire w_1738_;
wire w_1739_;
wire w_1740_;
wire w_1741_;
wire w_1742_;
wire w_1743_;
wire w_1744_;
wire w_1745_;
wire w_1746_;
wire w_1747_;
wire w_1748_;
wire w_1749_;
wire w_1750_;
wire w_1751_;
wire w_1752_;
wire w_1753_;
wire w_1754_;
wire w_1755_;
wire w_1756_;
wire w_1757_;
wire w_1758_;
wire w_1759_;
wire w_1760_;
wire w_1761_;
wire w_1762_;
wire w_1763_;
wire w_1764_;
wire w_1765_;
wire w_1766_;
wire w_1767_;
wire w_1768_;
wire w_1769_;
wire w_1770_;
wire w_1771_;
wire w_1772_;
wire w_1773_;
wire w_1774_;
wire w_1775_;
wire w_1776_;
wire w_1777_;
wire w_1778_;
wire w_1779_;
wire w_1780_;
wire w_1781_;
wire w_1782_;
wire w_1783_;
wire w_1784_;
wire w_1785_;
wire w_1786_;
wire w_1787_;
wire w_1788_;
wire w_1789_;
wire w_1790_;
wire w_1791_;
wire w_1792_;
wire w_1793_;
wire w_1794_;
wire w_1795_;
wire w_1796_;
wire w_1797_;
wire w_1798_;
wire w_1799_;
wire w_1800_;
wire w_1801_;
wire w_1802_;
wire w_1803_;
wire w_1804_;
wire w_1805_;
wire w_1806_;
wire w_1807_;
wire w_1808_;
wire w_1809_;
wire w_1810_;
wire w_1811_;
wire w_1812_;
wire w_1813_;
wire w_1814_;
wire w_1815_;
wire w_1816_;
wire w_1817_;
wire w_1818_;
wire w_1819_;
wire w_1820_;
wire w_1821_;
wire w_1822_;
wire w_1823_;
wire w_1824_;
wire w_1825_;
wire w_1826_;
wire w_1827_;
wire w_1828_;
wire w_1829_;
wire w_1830_;
wire w_1831_;
wire w_1832_;
wire w_1833_;
wire w_1834_;
wire w_1835_;
wire w_1836_;
wire w_1837_;
wire w_1838_;
wire w_1839_;
wire w_1840_;
wire w_1841_;
wire w_1842_;
wire w_1843_;
wire w_1844_;
wire w_1845_;
wire w_1846_;
wire w_1847_;
wire w_1848_;
wire w_1849_;
wire w_1850_;
wire w_1851_;
wire w_1852_;
wire w_1853_;
wire w_1854_;
wire w_1855_;
wire w_1856_;
wire w_1857_;
wire w_1858_;
wire w_1859_;
wire w_1860_;
wire w_1861_;
wire w_1862_;
wire w_1863_;
wire w_1864_;
wire w_1865_;
wire w_1866_;
wire w_1867_;
wire w_1868_;
wire w_1869_;
wire w_1870_;
wire w_1871_;
wire w_1872_;
wire w_1873_;
wire w_1874_;
wire w_1875_;
wire w_1876_;
wire w_1877_;
wire w_1878_;
wire w_1879_;
wire w_1880_;
wire w_1881_;
wire w_1882_;
wire w_1883_;
wire w_1884_;
wire w_1885_;
wire w_1886_;
wire w_1887_;
wire w_1888_;
wire w_1889_;
wire w_1890_;
wire w_1891_;
wire w_1892_;
wire w_1893_;
wire w_1894_;
wire w_1895_;
wire w_1896_;
wire w_1897_;
wire w_1898_;
wire w_1899_;
wire w_1900_;
wire w_1901_;
wire w_1902_;
wire w_1903_;
wire w_1904_;
wire w_1905_;
wire w_1906_;
wire w_1907_;
wire w_1908_;
wire w_1909_;
wire w_1910_;
wire w_1911_;
wire w_1912_;
wire w_1913_;
wire w_1914_;
wire w_1915_;
wire w_1916_;
wire w_1917_;
wire w_1918_;
wire w_1919_;
wire w_1920_;
wire w_1921_;
wire w_1922_;
wire w_1923_;
wire w_1924_;
wire w_1925_;
wire w_1926_;
wire w_1927_;
wire w_1928_;
wire w_1929_;
wire w_1930_;
wire w_1931_;
wire w_1932_;
wire w_1933_;
wire w_1934_;
wire w_1935_;
wire w_1936_;
wire w_1937_;
wire w_1938_;
wire w_1939_;
wire w_1940_;
wire w_1941_;
wire w_1942_;
wire w_1943_;
wire w_1944_;
wire w_1945_;
wire w_1946_;
wire w_1947_;
wire w_1948_;
wire w_1949_;
wire w_1950_;
wire w_1951_;
wire w_1952_;
wire w_1953_;
wire w_1954_;
wire w_1955_;
wire w_1956_;
wire w_1957_;
wire w_1958_;
wire w_1959_;
wire w_1960_;
wire w_1961_;
wire w_1962_;
wire w_1963_;
wire w_1964_;
wire w_1965_;
wire w_1966_;
wire w_1967_;
wire w_1968_;
wire w_1969_;
wire w_1970_;
wire w_1971_;
wire w_1972_;
wire w_1973_;
wire w_1974_;
wire w_1975_;
wire w_1976_;
wire w_1977_;
wire w_1978_;
wire w_1979_;
wire w_1980_;
wire w_1981_;
wire w_1982_;
wire w_1983_;
wire w_1984_;
wire w_1985_;
wire w_1986_;
wire w_1987_;
wire w_1988_;
wire w_1989_;
wire w_1990_;
wire w_1991_;
wire w_1992_;
wire w_1993_;
wire w_1994_;
wire w_1995_;
wire w_1996_;
wire w_1997_;
wire w_1998_;
wire w_1999_;
wire w_2000_;
wire w_2001_;
wire w_2002_;
wire w_2003_;
wire w_2004_;
wire w_2005_;
wire w_2006_;
wire w_2007_;
wire w_2008_;
wire w_2009_;
wire w_2010_;
wire w_2011_;
wire w_2012_;
wire w_2013_;
wire w_2014_;
wire w_2015_;
wire w_2016_;
wire w_2017_;
wire w_2018_;
wire w_2019_;
wire w_2020_;
wire w_2021_;
wire w_2022_;
wire w_2023_;
wire w_2024_;
wire w_2025_;
wire w_2026_;
wire w_2027_;
wire w_2028_;
wire w_2029_;
wire w_2030_;
wire w_2031_;
wire w_2032_;
wire w_2033_;
wire w_2034_;
wire w_2035_;
wire w_2036_;
wire w_2037_;
wire w_2038_;
wire w_2039_;
wire w_2040_;
wire w_2041_;
wire w_2042_;
wire w_2043_;
wire w_2044_;
wire w_2045_;
wire w_2046_;
wire w_2047_;
wire w_2048_;
wire w_2049_;
wire w_2050_;
wire w_2051_;
wire w_2052_;
wire w_2053_;
wire w_2054_;
wire w_2055_;
wire w_2056_;
wire w_2057_;
wire w_2058_;
wire w_2059_;
wire w_2060_;
wire w_2061_;
wire w_2062_;
wire w_2063_;
wire w_2064_;
wire w_2065_;
wire w_2066_;
wire w_2067_;
wire w_2068_;
wire w_2069_;
wire w_2070_;
wire w_2071_;
wire w_2072_;
wire w_2073_;
wire w_2074_;
wire w_2075_;
wire w_2076_;
wire w_2077_;
wire w_2078_;
wire w_2079_;
wire w_2080_;
wire w_2081_;
wire w_2082_;
wire w_2083_;
wire w_2084_;
wire w_2085_;
wire w_2086_;
wire w_2087_;
wire w_2088_;
wire w_2089_;
wire w_2090_;
wire w_2091_;
wire w_2092_;
wire w_2093_;
wire w_2094_;
wire w_2095_;
wire w_2096_;
wire w_2097_;
wire w_2098_;
wire w_2099_;
wire w_2100_;
wire w_2101_;
wire w_2102_;
wire w_2103_;
wire w_2104_;
wire w_2105_;
wire w_2106_;
wire w_2107_;
wire w_2108_;
wire w_2109_;
wire w_2110_;
wire w_2111_;
wire w_2112_;
wire w_2113_;
wire w_2114_;
wire w_2115_;
wire w_2116_;
wire w_2117_;
wire w_2118_;
wire w_2119_;
wire w_2120_;
wire w_2121_;
wire w_2122_;
wire w_2123_;
wire w_2124_;
wire w_2125_;
wire w_2126_;
wire w_2127_;
wire w_2128_;
wire w_2129_;
wire w_2130_;
wire w_2131_;
wire w_2132_;
wire w_2133_;
wire w_2134_;
wire w_2135_;
wire w_2136_;
wire w_2137_;
wire w_2138_;
wire w_2139_;
wire w_2140_;
wire w_2141_;
wire w_2142_;
wire w_2143_;
wire w_2144_;
wire w_2145_;
wire w_2146_;
wire w_2147_;
wire w_2148_;
wire w_2149_;
wire w_2150_;
wire w_2151_;
wire w_2152_;
wire w_2153_;
wire w_2154_;
wire w_2155_;
wire w_2156_;
wire w_2157_;
wire w_2158_;
wire w_2159_;
wire w_2160_;
wire w_2161_;
wire w_2162_;
wire w_2163_;
wire w_2164_;
wire w_2165_;
wire w_2166_;
wire w_2167_;
wire w_2168_;
wire w_2169_;
wire w_2170_;
wire w_2171_;
wire w_2172_;
wire w_2173_;
wire w_2174_;
wire w_2175_;
wire w_2176_;
wire w_2177_;
wire w_2178_;
wire w_2179_;
wire w_2180_;
wire w_2181_;
wire w_2182_;
wire w_2183_;
wire w_2184_;
wire w_2185_;
wire w_2186_;
wire w_2187_;
wire w_2188_;
wire w_2189_;
wire w_2190_;
wire w_2191_;
wire w_2192_;
wire w_2193_;
wire w_2194_;
wire w_2195_;
wire w_2196_;
wire w_2197_;
wire w_2198_;
wire w_2199_;
wire w_2200_;
wire w_2201_;
wire w_2202_;
wire w_2203_;
wire w_2204_;
wire w_2205_;
wire w_2206_;
wire w_2207_;
wire w_2208_;
wire w_2209_;
wire w_2210_;
wire w_2211_;
wire w_2212_;
wire w_2213_;
wire w_2214_;
wire w_2215_;
wire w_2216_;
wire w_2217_;
wire w_2218_;
wire w_2219_;
wire w_2220_;
wire w_2221_;
wire w_2222_;
wire w_2223_;
wire w_2224_;
wire w_2225_;
wire w_2226_;
wire w_2227_;
wire w_2228_;
wire w_2229_;
wire w_2230_;
wire w_2231_;
wire w_2232_;
wire w_2233_;
wire w_2234_;
wire w_2235_;
wire w_2236_;
wire w_2237_;
wire w_2238_;
wire w_2239_;
wire w_2240_;
wire w_2241_;
wire w_2242_;
wire w_2243_;
wire w_2244_;
wire w_2245_;
wire w_2246_;
wire w_2247_;
wire w_2248_;
wire w_2249_;
wire w_2250_;
wire w_2251_;
wire w_2252_;
wire w_2253_;
wire w_2254_;
wire w_2255_;
wire w_2256_;
wire w_2257_;
wire w_2258_;
wire w_2259_;
wire w_2260_;
wire w_2261_;
wire w_2262_;
wire w_2263_;
wire w_2264_;
wire w_2265_;
wire w_2266_;
wire w_2267_;
wire w_2268_;
wire w_2269_;
wire w_2270_;
wire w_2271_;
wire w_2272_;
wire w_2273_;
wire w_2274_;
wire w_2275_;
wire w_2276_;
wire w_2277_;
wire w_2278_;
wire w_2279_;
wire w_2280_;
wire w_2281_;
wire w_2282_;
wire w_2283_;
wire w_2284_;
wire w_2285_;
wire w_2286_;
wire w_2287_;
wire w_2288_;
wire w_2289_;
wire w_2290_;
wire w_2291_;
wire w_2292_;
wire w_2293_;
wire w_2294_;
wire w_2295_;
wire w_2296_;
wire w_2297_;
wire w_2298_;
wire w_2299_;
wire w_2300_;
wire w_2301_;
wire w_2302_;
wire w_2303_;
wire w_2304_;
wire w_2305_;
wire w_2306_;
wire w_2307_;
wire w_2308_;
wire w_2309_;
wire w_2310_;
wire w_2311_;
wire w_2312_;
wire w_2313_;
wire w_2314_;
wire w_2315_;
wire w_2316_;
wire w_2317_;
wire w_2318_;
wire w_2319_;
wire w_2320_;
wire w_2321_;
wire w_2322_;
wire w_2323_;
wire w_2324_;
wire w_2325_;
wire w_2326_;
wire w_2327_;
wire w_2328_;
wire w_2329_;
wire w_2330_;
wire w_2331_;
wire w_2332_;
wire w_2333_;
wire w_2334_;
wire w_2335_;
wire w_2336_;
wire w_2337_;
wire w_2338_;
wire w_2339_;
wire w_2340_;
wire w_2341_;
wire w_2342_;
wire w_2343_;
wire w_2344_;
wire w_2345_;
wire w_2346_;
wire w_2347_;
wire w_2348_;
wire w_2349_;
wire w_2350_;
wire w_2351_;
wire w_2352_;
wire w_2353_;
wire w_2354_;
wire w_2355_;
wire w_2356_;
wire w_2357_;
wire w_2358_;
wire w_2359_;
wire w_2360_;
wire w_2361_;
wire w_2362_;
wire w_2363_;
wire w_2364_;
wire w_2365_;
wire w_2366_;
wire w_2367_;
wire w_2368_;
wire w_2369_;
wire w_2370_;
wire w_2371_;
wire w_2372_;
wire w_2373_;
wire w_2374_;
wire w_2375_;
wire w_2376_;
wire w_2377_;
wire w_2378_;
wire w_2379_;
wire w_2380_;
wire w_2381_;
wire w_2382_;
wire w_2383_;
wire w_2384_;
wire w_2385_;
wire w_2386_;
wire w_2387_;
wire w_2388_;
wire w_2389_;
wire w_2390_;
wire w_2391_;
wire w_2392_;
wire w_2393_;
wire w_2394_;
wire w_2395_;
wire w_2396_;
wire w_2397_;
wire w_2398_;
wire w_2399_;
wire w_2400_;
wire w_2401_;
wire w_2402_;
wire w_2403_;
wire w_2404_;
wire w_2405_;
wire w_2406_;
wire w_2407_;
wire w_2408_;
wire w_2409_;
wire w_2410_;
wire w_2411_;
wire w_2412_;
wire w_2413_;
wire w_2414_;
wire w_2415_;
wire w_2416_;
wire w_2417_;
wire w_2418_;
wire w_2419_;
wire w_2420_;
wire w_2421_;
wire w_2422_;
wire w_2423_;
wire w_2424_;
wire w_2425_;
wire w_2426_;
wire w_2427_;
wire w_2428_;
wire w_2429_;
wire w_2430_;
wire w_2431_;
wire w_2432_;
wire w_2433_;
wire w_2434_;
wire w_2435_;
wire w_2436_;
wire w_2437_;
wire w_2438_;
wire w_2439_;
wire w_2440_;
wire w_2441_;
wire w_2442_;
wire w_2443_;
wire w_2444_;
wire w_2445_;
wire w_2446_;
wire w_2447_;
wire w_2448_;
wire w_2449_;
wire w_2450_;
wire w_2451_;
wire w_2452_;
wire w_2453_;
wire w_2454_;
wire w_2455_;
wire w_2456_;
wire w_2457_;
wire w_2458_;
wire w_2459_;
wire w_2460_;
wire w_2461_;
wire w_2462_;
wire w_2463_;
wire w_2464_;
wire w_2465_;
wire w_2466_;
wire w_2467_;
wire w_2468_;
wire w_2469_;
wire w_2470_;
wire w_2471_;
wire w_2472_;
wire w_2473_;
wire w_2474_;
wire w_2475_;
wire w_2476_;
wire w_2477_;
wire w_2478_;
wire w_2479_;
wire w_2480_;
wire w_2481_;
wire w_2482_;
wire w_2483_;
wire w_2484_;
wire w_2485_;
wire w_2486_;
wire w_2487_;
wire w_2488_;
wire w_2489_;
wire w_2490_;
wire w_2491_;
wire w_2492_;
wire w_2493_;
wire w_2494_;
wire w_2495_;
wire w_2496_;
wire w_2497_;
wire w_2498_;
wire w_2499_;
wire w_2500_;
wire w_2501_;
wire w_2502_;
wire w_2503_;
wire w_2504_;
wire w_2505_;
wire w_2506_;
wire w_2507_;
wire w_2508_;
wire w_2509_;
wire w_2510_;
wire w_2511_;
wire w_2512_;
wire w_2513_;
wire w_2514_;
wire w_2515_;
wire w_2516_;
wire w_2517_;
wire w_2518_;
wire w_2519_;
wire w_2520_;
wire w_2521_;
wire w_2522_;
wire w_2523_;
wire w_2524_;
wire w_2525_;
wire w_2526_;
wire w_2527_;
wire w_2528_;
wire w_2529_;
wire w_2530_;
wire w_2531_;
wire w_2532_;
wire w_2533_;
wire w_2534_;
wire w_2535_;
wire w_2536_;
wire w_2537_;
wire w_2538_;
wire w_2539_;
wire w_2540_;
wire w_2541_;
wire w_2542_;
wire w_2543_;
wire w_2544_;
wire w_2545_;
wire w_2546_;
wire w_2547_;
wire w_2548_;
wire w_2549_;
wire w_2550_;
wire w_2551_;
wire w_2552_;
wire w_2553_;
wire w_2554_;
wire w_2555_;
wire w_2556_;
wire w_2557_;
wire w_2558_;
wire w_2559_;
wire w_2560_;
wire w_2561_;
wire w_2562_;
wire w_2563_;
wire w_2564_;
wire w_2565_;
wire w_2566_;
wire w_2567_;
wire w_2568_;
wire w_2569_;
wire w_2570_;
wire w_2571_;
wire w_2572_;
wire w_2573_;
wire w_2574_;
wire w_2575_;
wire w_2576_;
wire w_2577_;
wire w_2578_;
wire w_2579_;
wire w_2580_;
wire w_2581_;
wire w_2582_;
wire w_2583_;
wire w_2584_;
wire w_2585_;
wire w_2586_;
wire w_2587_;
wire w_2588_;
wire w_2589_;
wire w_2590_;
wire w_2591_;
wire w_2592_;
wire w_2593_;
wire w_2594_;
wire w_2595_;
wire w_2596_;
wire w_2597_;
wire w_2598_;
wire w_2599_;
wire w_2600_;
wire w_2601_;
wire w_2602_;
wire w_2603_;
wire w_2604_;
wire w_2605_;
wire w_2606_;
wire w_2607_;
wire w_2608_;
wire w_2609_;
wire w_2610_;
wire w_2611_;
wire w_2612_;
wire w_2613_;
wire w_2614_;
wire w_2615_;
wire w_2616_;
wire w_2617_;
wire w_2618_;
wire w_2619_;
wire w_2620_;
wire w_2621_;
wire w_2622_;
wire w_2623_;
wire w_2624_;
wire w_2625_;
wire w_2626_;
wire w_2627_;
wire w_2628_;
wire w_2629_;
wire w_2630_;
wire w_2631_;
wire w_2632_;
wire w_2633_;
wire w_2634_;
wire w_2635_;
wire w_2636_;
wire w_2637_;
wire w_2638_;
wire w_2639_;
wire w_2640_;
wire w_2641_;
wire w_2642_;
wire w_2643_;
wire w_2644_;
wire w_2645_;
wire w_2646_;
wire w_2647_;
wire w_2648_;
wire w_2649_;
wire w_2650_;
wire w_2651_;
wire w_2652_;
wire w_2653_;
wire w_2654_;
wire w_2655_;
wire w_2656_;
wire w_2657_;
wire w_2658_;
wire w_2659_;
wire w_2660_;
wire w_2661_;
wire w_2662_;
wire w_2663_;
wire w_2664_;
wire w_2665_;
wire w_2666_;
wire w_2667_;
wire w_2668_;
wire w_2669_;
wire w_2670_;
wire w_2671_;
wire w_2672_;
wire w_2673_;
wire w_2674_;
wire w_2675_;
wire w_2676_;
wire w_2677_;
wire w_2678_;
wire w_2679_;
wire w_2680_;
wire w_2681_;
wire w_2682_;
wire w_2683_;
wire w_2684_;
wire w_2685_;
wire w_2686_;
wire w_2687_;
wire w_2688_;
wire w_2689_;
wire w_2690_;
wire w_2691_;
wire w_2692_;
wire w_2693_;
wire w_2694_;
wire w_2695_;
wire w_2696_;
wire w_2697_;
wire w_2698_;
wire w_2699_;
wire w_2700_;
wire w_2701_;
wire w_2702_;
wire w_2703_;
wire w_2704_;
wire w_2705_;
wire w_2706_;
wire w_2707_;
wire w_2708_;
wire w_2709_;
wire w_2710_;
wire w_2711_;
wire w_2712_;
wire w_2713_;
wire w_2714_;
wire w_2715_;
wire w_2716_;
wire w_2717_;
wire w_2718_;
wire w_2719_;
wire w_2720_;
wire w_2721_;
wire w_2722_;
wire w_2723_;
wire w_2724_;
wire w_2725_;
wire w_2726_;
wire w_2727_;
wire w_2728_;
wire w_2729_;
wire w_2730_;
wire w_2731_;
wire w_2732_;
wire w_2733_;
wire w_2734_;
wire w_2735_;
wire w_2736_;
wire w_2737_;
wire w_2738_;
wire w_2739_;
wire w_2740_;
wire w_2741_;
wire w_2742_;
wire w_2743_;
wire w_2744_;
wire w_2745_;
wire w_2746_;
wire w_2747_;
wire w_2748_;
wire w_2749_;
wire w_2750_;
wire w_2751_;
wire w_2752_;
wire w_2753_;
wire w_2754_;
wire w_2755_;
wire w_2756_;
wire w_2757_;
wire w_2758_;
wire w_2759_;
wire w_2760_;
wire w_2761_;
wire w_2762_;
wire w_2763_;
wire w_2764_;
wire w_2765_;
wire w_2766_;
wire w_2767_;
wire w_2768_;
wire w_2769_;
wire w_2770_;
wire w_2771_;
wire w_2772_;
wire w_2773_;
wire w_2774_;
wire w_2775_;
wire w_2776_;
wire w_2777_;
wire w_2778_;
wire w_2779_;
wire w_2780_;
wire w_2781_;
wire w_2782_;
wire w_2783_;
wire w_2784_;
wire w_2785_;
wire w_2786_;
wire w_2787_;
wire w_2788_;
wire w_2789_;
wire w_2790_;
wire w_2791_;
wire w_2792_;
wire w_2793_;
wire w_2794_;
wire w_2795_;
wire w_2796_;
wire w_2797_;
wire w_2798_;
wire w_2799_;
wire w_2800_;
wire w_2801_;
wire w_2802_;
wire w_2803_;
wire w_2804_;
wire w_2805_;
wire w_2806_;
wire w_2807_;
wire w_2808_;
wire w_2809_;
wire w_2810_;
wire w_2811_;
wire w_2812_;
wire w_2813_;
wire w_2814_;
wire w_2815_;
wire w_2816_;
wire w_2817_;
wire w_2818_;
wire w_2819_;
wire w_2820_;
wire w_2821_;
wire w_2822_;
wire w_2823_;
wire w_2824_;
wire w_2825_;
wire w_2826_;
wire w_2827_;
wire w_2828_;
wire w_2829_;
wire w_2830_;
wire w_2831_;
wire w_2832_;
wire w_2833_;
wire w_2834_;
wire w_2835_;
wire w_2836_;
wire w_2837_;
wire w_2838_;
wire w_2839_;
wire w_2840_;
wire w_2841_;
wire w_2842_;
wire w_2843_;
wire w_2844_;
wire w_2845_;
wire w_2846_;
wire w_2847_;
wire w_2848_;
wire w_2849_;
wire w_2850_;
wire w_2851_;
wire w_2852_;
wire w_2853_;
wire w_2854_;
wire w_2855_;
wire w_2856_;
wire w_2857_;
wire w_2858_;
wire w_2859_;
wire w_2860_;
wire w_2861_;
wire w_2862_;
wire w_2863_;
wire w_2864_;
wire w_2865_;
wire w_2866_;
wire w_2867_;
wire w_2868_;
wire w_2869_;
wire w_2870_;
wire w_2871_;
wire w_2872_;
wire w_2873_;
wire w_2874_;
wire w_2875_;
wire w_2876_;
wire w_2877_;
wire w_2878_;
wire w_2879_;
wire w_2880_;
wire w_2881_;
wire w_2882_;
wire w_2883_;
wire w_2884_;
wire w_2885_;
wire w_2886_;
wire w_2887_;
wire w_2888_;
wire w_2889_;
wire w_2890_;
wire w_2891_;
wire w_2892_;
wire w_2893_;
wire w_2894_;
wire w_2895_;
wire w_2896_;
wire w_2897_;
wire w_2898_;
wire w_2899_;
wire w_2900_;
wire w_2901_;
wire w_2902_;
wire w_2903_;
wire w_2904_;
wire w_2905_;
wire w_2906_;
wire w_2907_;
wire w_2908_;
wire w_2909_;
wire w_2910_;
wire w_2911_;
wire w_2912_;
wire w_2913_;
wire w_2914_;
wire w_2915_;
wire w_2916_;
wire w_2917_;
wire w_2918_;
wire w_2919_;
wire w_2920_;
wire w_2921_;
wire w_2922_;
wire w_2923_;
wire w_2924_;
wire w_2925_;
wire w_2926_;
wire w_2927_;
wire w_2928_;
wire w_2929_;
wire w_2930_;
wire w_2931_;
wire w_2932_;
wire w_2933_;
wire w_2934_;
wire w_2935_;
wire w_2936_;
wire w_2937_;
wire w_2938_;
wire w_2939_;
wire w_2940_;
wire w_2941_;
wire w_2942_;
wire w_2943_;
wire w_2944_;
wire w_2945_;
wire w_2946_;
wire w_2947_;
wire w_2948_;
wire w_2949_;
wire w_2950_;
wire w_2951_;
wire w_2952_;
wire w_2953_;
wire w_2954_;
wire w_2955_;
wire w_2956_;
wire w_2957_;
wire w_2958_;
wire w_2959_;
wire w_2960_;
wire w_2961_;
wire w_2962_;
wire w_2963_;
wire w_2964_;
wire w_2965_;
wire w_2966_;
wire w_2967_;
wire w_2968_;
wire w_2969_;
wire w_2970_;
wire w_2971_;
wire w_2972_;
wire w_2973_;
wire w_2974_;
wire w_2975_;
wire w_2976_;
wire w_2977_;
wire w_2978_;
wire w_2979_;
wire w_2980_;
wire w_2981_;
wire w_2982_;
wire w_2983_;
wire w_2984_;
wire w_2985_;
wire w_2986_;
wire w_2987_;
wire w_2988_;
wire w_2989_;
wire w_2990_;
wire w_2991_;
wire w_2992_;
wire w_2993_;
wire w_2994_;
wire w_2995_;
wire w_2996_;
wire w_2997_;
wire w_2998_;
wire w_2999_;
wire w_3000_;
wire w_3001_;
wire w_3002_;
wire w_3003_;
wire w_3004_;
wire w_3005_;
wire w_3006_;
wire w_3007_;
wire w_3008_;
wire w_3009_;
wire w_3010_;
wire w_3011_;
wire w_3012_;
wire w_3013_;
wire w_3014_;
wire w_3015_;
wire w_3016_;
wire w_3017_;
wire w_3018_;
wire w_3019_;
wire w_3020_;
wire w_3021_;
wire w_3022_;
wire w_3023_;
wire w_3024_;
wire w_3025_;
wire w_3026_;
wire w_3027_;
wire w_3028_;
wire w_3029_;
wire w_3030_;
wire w_3031_;
wire w_3032_;
wire w_3033_;
wire w_3034_;
wire w_3035_;
wire w_3036_;
wire w_3037_;
wire w_3038_;
wire w_3039_;
wire w_3040_;
wire w_3041_;
wire w_3042_;
wire w_3043_;
wire w_3044_;
wire w_3045_;
wire w_3046_;
wire w_3047_;
wire w_3048_;
wire w_3049_;
wire w_3050_;
wire w_3051_;
wire w_3052_;
wire w_3053_;
wire w_3054_;
wire w_3055_;
wire w_3056_;
wire w_3057_;
wire w_3058_;
wire w_3059_;
wire w_3060_;
wire w_3061_;
wire w_3062_;
wire w_3063_;
wire w_3064_;
wire w_3065_;
wire w_3066_;
wire w_3067_;
wire w_3068_;
wire w_3069_;
wire w_3070_;
wire w_3071_;
wire w_3072_;
wire w_3073_;
wire w_3074_;
wire w_3075_;
wire w_3076_;
wire w_3077_;
wire w_3078_;
wire w_3079_;
wire w_3080_;
wire w_3081_;
wire w_3082_;
wire w_3083_;
wire w_3084_;
wire w_3085_;
wire w_3086_;
wire w_3087_;
wire w_3088_;
wire w_3089_;
wire w_3090_;
wire w_3091_;
wire w_3092_;
wire w_3093_;
wire w_3094_;
wire w_3095_;
wire w_3096_;
wire w_3097_;
wire w_3098_;
wire w_3099_;
wire w_3100_;
wire w_3101_;
wire w_3102_;
wire w_3103_;
wire w_3104_;
wire w_3105_;
wire w_3106_;
wire w_3107_;
wire w_3108_;
wire w_3109_;
wire w_3110_;
wire w_3111_;
wire w_3112_;
wire w_3113_;
wire w_3114_;
wire w_3115_;
wire w_3116_;
wire w_3117_;
wire w_3118_;
wire w_3119_;
wire w_3120_;
wire w_3121_;
wire w_3122_;
wire w_3123_;
wire w_3124_;
wire w_3125_;
wire w_3126_;
wire w_3127_;
wire w_3128_;
wire w_3129_;
wire w_3130_;
wire w_3131_;
wire w_3132_;
wire w_3133_;
wire w_3134_;
wire w_3135_;
wire w_3136_;
wire w_3137_;
wire w_3138_;
wire w_3139_;
wire w_3140_;
wire w_3141_;
wire w_3142_;
wire w_3143_;
wire w_3144_;
wire w_3145_;
wire w_3146_;
wire w_3147_;
wire w_3148_;
wire w_3149_;
wire w_3150_;
wire w_3151_;
wire w_3152_;
wire w_3153_;
wire w_3154_;
wire w_3155_;
wire w_3156_;
wire w_3157_;
wire w_3158_;
wire w_3159_;
wire w_3160_;
wire w_3161_;
wire w_3162_;
wire w_3163_;
wire w_3164_;
wire w_3165_;
wire w_3166_;
wire w_3167_;
wire w_3168_;
wire w_3169_;
wire w_3170_;
wire w_3171_;
wire w_3172_;
wire w_3173_;
wire w_3174_;
wire w_3175_;
wire w_3176_;
wire w_3177_;
wire w_3178_;
wire w_3179_;
wire w_3180_;
wire w_3181_;
wire w_3182_;
wire w_3183_;
wire w_3184_;
wire w_3185_;
wire w_3186_;
wire w_3187_;
wire w_3188_;
wire w_3189_;
wire w_3190_;
wire w_3191_;
wire w_3192_;
wire w_3193_;
wire w_3194_;
wire w_3195_;
wire w_3196_;
wire w_3197_;
wire w_3198_;
wire w_3199_;
wire w_3200_;
wire w_3201_;
wire w_3202_;
wire w_3203_;
wire w_3204_;
wire w_3205_;
wire w_3206_;
wire w_3207_;
wire w_3208_;
wire w_3209_;
wire w_3210_;
wire w_3211_;
wire w_3212_;
wire w_3213_;
wire w_3214_;
wire w_3215_;
wire w_3216_;
wire w_3217_;
wire w_3218_;
wire w_3219_;
wire w_3220_;
wire w_3221_;
wire w_3222_;
wire w_3223_;
wire w_3224_;
wire w_3225_;
wire w_3226_;
wire w_3227_;
wire w_3228_;
wire w_3229_;
wire w_3230_;
wire w_3231_;
wire w_3232_;
wire w_3233_;
wire w_3234_;
wire w_3235_;
wire w_3236_;
wire w_3237_;
wire w_3238_;
wire w_3239_;
wire w_3240_;
wire w_3241_;
wire w_3242_;
wire w_3243_;
wire w_3244_;
wire w_3245_;
wire w_3246_;
wire w_3247_;
wire w_3248_;
wire w_3249_;
wire w_3250_;
wire w_3251_;
wire w_3252_;
wire w_3253_;
wire w_3254_;
wire w_3255_;
wire w_3256_;
wire w_3257_;
wire w_3258_;
wire w_3259_;
wire w_3260_;
wire w_3261_;
wire w_3262_;
wire w_3263_;
wire w_3264_;
wire w_3265_;
wire w_3266_;
wire w_3267_;
wire w_3268_;
wire w_3269_;
wire w_3270_;
wire w_3271_;
wire w_3272_;
wire w_3273_;
wire w_3274_;
wire w_3275_;
wire w_3276_;
wire w_3277_;
wire w_3278_;
wire w_3279_;
wire w_3280_;
wire w_3281_;
wire w_3282_;
wire w_3283_;
wire w_3284_;
wire w_3285_;
wire w_3286_;
wire w_3287_;
wire w_3288_;
wire w_3289_;
wire w_3290_;
wire w_3291_;
wire w_3292_;
wire w_3293_;
wire w_3294_;
wire w_3295_;
wire w_3296_;
wire w_3297_;
wire w_3298_;
wire w_3299_;
wire w_3300_;
wire w_3301_;
wire w_3302_;
wire w_3303_;
wire w_3304_;
wire w_3305_;
wire w_3306_;
wire w_3307_;
wire w_3308_;
wire w_3309_;
wire w_3310_;
wire w_3311_;
wire w_3312_;
wire w_3313_;
wire w_3314_;
wire w_3315_;
wire w_3316_;
wire w_3317_;
wire w_3318_;
wire w_3319_;
wire w_3320_;
wire w_3321_;
wire w_3322_;
wire w_3323_;
wire w_3324_;
wire w_3325_;
wire w_3326_;
wire w_3327_;
wire w_3328_;
wire w_3329_;
wire w_3330_;
wire w_3331_;
wire w_3332_;
wire w_3333_;
wire w_3334_;
wire w_3335_;
wire w_3336_;
wire w_3337_;
wire w_3338_;
wire w_3339_;
wire w_3340_;
wire w_3341_;
wire w_3342_;
wire w_3343_;
wire w_3344_;
wire w_3345_;
wire w_3346_;
wire w_3347_;
wire w_3348_;
wire w_3349_;
wire w_3350_;
wire w_3351_;
wire w_3352_;
wire w_3353_;
wire w_3354_;
wire w_3355_;
wire w_3356_;
wire w_3357_;
wire w_3358_;
wire w_3359_;
wire w_3360_;
wire w_3361_;
wire w_3362_;
wire w_3363_;
wire w_3364_;
wire w_3365_;
wire w_3366_;
wire w_3367_;
wire w_3368_;
wire w_3369_;
wire w_3370_;
wire w_3371_;
wire w_3372_;
wire w_3373_;
wire w_3374_;
wire w_3375_;
wire w_3376_;
wire w_3377_;
wire w_3378_;
wire w_3379_;
wire w_3380_;
wire w_3381_;
wire w_3382_;
wire w_3383_;
wire w_3384_;
wire w_3385_;
wire w_3386_;
wire w_3387_;
wire w_3388_;
wire w_3389_;
wire w_3390_;
wire w_3391_;
wire w_3392_;
wire w_3393_;
wire w_3394_;
wire w_3395_;
wire w_3396_;
wire w_3397_;
wire w_3398_;
wire w_3399_;
wire w_3400_;
wire w_3401_;
wire w_3402_;
wire w_3403_;
wire w_3404_;
wire w_3405_;
wire w_3406_;
wire w_3407_;
wire w_3408_;
wire w_3409_;
wire w_3410_;
wire w_3411_;
wire w_3412_;
wire w_3413_;
wire w_3414_;
wire w_3415_;
wire w_3416_;
wire w_3417_;
wire w_3418_;
wire w_3419_;
wire w_3420_;
wire w_3421_;
wire w_3422_;
wire w_3423_;
wire w_3424_;
wire w_3425_;
wire w_3426_;
wire w_3427_;
wire w_3428_;
wire w_3429_;
wire w_3430_;
wire w_3431_;
wire w_3432_;
wire w_3433_;
wire w_3434_;
wire w_3435_;
wire w_3436_;
wire w_3437_;
wire w_3438_;
wire w_3439_;
wire w_3440_;
wire w_3441_;
wire w_3442_;
wire w_3443_;
wire w_3444_;
wire w_3445_;
wire w_3446_;
wire w_3447_;
wire w_3448_;
wire w_3449_;
wire w_3450_;
wire w_3451_;
wire w_3452_;
wire w_3453_;
wire w_3454_;
wire w_3455_;
wire w_3456_;
wire w_3457_;
wire w_3458_;
wire w_3459_;
wire w_3460_;
wire w_3461_;
wire w_3462_;
wire w_3463_;
wire w_3464_;
wire w_3465_;
wire w_3466_;
wire w_3467_;
wire w_3468_;
wire w_3469_;
wire w_3470_;
wire w_3471_;
wire w_3472_;
wire w_3473_;
wire w_3474_;
wire w_3475_;
wire w_3476_;
wire w_3477_;
wire w_3478_;
wire w_3479_;
wire w_3480_;
wire w_3481_;
wire w_3482_;
wire w_3483_;
wire w_3484_;
wire w_3485_;
wire w_3486_;
wire w_3487_;
wire w_3488_;
wire w_3489_;
wire w_3490_;
wire w_3491_;
wire w_3492_;
wire w_3493_;
wire w_3494_;
wire w_3495_;
wire w_3496_;
wire w_3497_;
wire w_3498_;
wire w_3499_;
wire w_3500_;
wire w_3501_;
wire w_3502_;
wire w_3503_;
wire w_3504_;
wire w_3505_;
wire w_3506_;
wire w_3507_;
wire w_3508_;
wire w_3509_;
wire w_3510_;
wire w_3511_;
wire w_3512_;
wire w_3513_;
wire w_3514_;
wire w_3515_;
wire w_3516_;
wire w_3517_;
wire w_3518_;
wire w_3519_;
wire w_3520_;
wire w_3521_;
wire w_3522_;
wire w_3523_;
wire w_3524_;
wire w_3525_;
wire w_3526_;
wire w_3527_;
wire w_3528_;
or (w_2367_, w_1842_, w_1474_);
or (w_0651_, in5[2], w_2063_);
and (w_0912_, w_0002_, w_2955_);
not (w_2710_, w_1297_);
or (w_1236_, w_2707_, w_1751_);
not (w_3267_, w_1141_);
and (w_1759_, w_2563_, w_0599_);
or (w_2551_, w_2263_, w_2391_);
not (w_0165_, in2[1]);
or (w_2977_, in7[4], w_2229_);
or (out8[3], w_1731_, w_0556_);
or (out18[7], w_2518_, w_1022_);
and (w_2982_, in14[7], w_2482_);
or (w_2593_, w_0680_, w_0055_);
and (out1[1], w_3067_, w_2930_);
or (w_3163_, w_0850_, w_1581_);
or (w_0998_, w_1240_, w_2824_);
and (w_2494_, w_3173_, w_1157_);
and (w_0188_, in9[1], in10[1]);
and (w_1743_, w_2397_, w_2682_);
or (out11[3], w_1077_, w_1652_);
or (w_1133_, w_2732_, w_2527_);
not (w_0385_, in10[0]);
and (w_2226_, in16[1], w_0208_);
or (w_3186_, w_2364_, w_2309_);
or (w_1938_, w_0781_, w_1683_);
and (w_1828_, in3[0], w_0328_);
not (w_2415_, w_0666_);
and (w_2567_, w_1616_, w_2545_);
not (w_0970_, in4[2]);
and (w_2848_, w_2305_, w_2298_);
or (w_2675_, w_2864_, w_1891_);
not (w_0543_, in5[2]);
and (w_2563_, w_2793_, w_1914_);
or (w_1214_, w_0416_, w_1989_);
or (out16[6], w_3349_, w_2008_);
and (w_1838_, w_2270_, w_0405_);
or (w_2690_, w_0970_, w_0902_);
not (w_2137_, in13[0]);
and (w_0295_, w_1423_, w_2464_);
or (w_2199_, w_2753_, w_2043_);
and (w_3191_, w_2827_, w_0066_);
or (out5[0], w_2326_, w_2951_);
and (w_2122_, w_0842_, w_1334_);
not (w_3500_, w_3115_);
or (w_1299_, w_2371_, w_1791_);
and (w_1052_, w_1202_, w_2332_);
and (w_3502_, w_3282_, w_1700_);
and (w_2048_, w_1541_, w_3162_);
or (w_3444_, w_2060_, w_1003_);
and (w_1282_, w_1025_, w_3343_);
or (w_1293_, in15[4], w_3026_);
not (w_3215_, in10[1]);
and (out24[4], w_0087_, w_1579_);
and (w_2324_, w_1291_, w_2070_);
and (w_1148_, w_1355_, w_2367_);
and (w_3225_, in6[3], w_3483_);
not (w_2742_, w_0331_);
and (w_2282_, w_3029_, w_2626_);
not (w_2256_, w_1833_);
and (w_0624_, w_0991_, w_1233_);
or (w_1889_, w_2650_, w_2680_);
or (w_2801_, w_1320_, w_2131_);
and (w_3359_, w_0992_, w_0003_);
and (w_0796_, in8[5], w_1076_);
and (w_0397_, w_1183_, w_2783_);
or (w_3307_, in1[2], in2[2]);
not (w_0767_, w_3055_);
or (w_2375_, in4[5], w_2945_);
or (out20[7], w_0168_, w_0357_);
and (w_1905_, w_1033_, w_0304_);
or (w_2374_, w_1274_, w_0404_);
not (w_0534_, w_2706_);
or (w_3004_, w_1014_, w_1231_);
or (w_3504_, w_0443_, w_0976_);
and (w_1627_, w_2563_, w_3021_);
or (w_0550_, w_2277_, w_2826_);
and (w_3247_, w_1876_, w_3183_);
and (w_3049_, w_2955_, w_2320_);
or (w_2731_, w_1320_, w_1714_);
and (w_1825_, w_0780_, w_0292_);
and (w_1141_, w_2134_, w_1785_);
or (w_2314_, w_2303_, w_2622_);
or (w_0944_, w_3446_, w_1812_);
or (w_3239_, w_2470_, w_2612_);
and (w_1667_, w_3048_, w_2102_);
and (w_3284_, w_0413_, w_1677_);
or (w_0252_, w_0136_, w_0491_);
or (w_1784_, w_3070_, w_0558_);
or (out9[3], w_1554_, w_0566_);
and (w_1461_, w_0013_, w_0845_);
and (w_1842_, w_2584_, w_3381_);
and (w_2637_, w_0629_, w_3118_);
and (w_0622_, in4[5], w_1922_);
or (w_0411_, in9[3], in10[3]);
not (w_2156_, w_1488_);
or (w_2821_, w_0322_, w_2778_);
or (w_1451_, in11[5], w_3479_);
not (w_0215_, in3[5]);
or (w_0074_, w_0365_, w_2275_);
or (w_1013_, w_0982_, w_3177_);
or (w_1319_, w_2694_, w_3190_);
and (w_3010_, w_1236_, w_3291_);
not (w_0373_, w_2215_);
or (w_1344_, w_2618_, w_2042_);
or (w_1843_, w_2460_, w_3016_);
and (w_1926_, w_2961_, w_1192_);
and (w_3169_, w_3445_, w_0650_);
or (w_3379_, w_0654_, w_3097_);
and (w_2327_, w_1243_, w_0881_);
and (w_2940_, w_0452_, w_0897_);
or (w_3305_, in12[3], w_1748_);
or (w_1541_, w_1655_, w_0448_);
or (w_2503_, w_2005_, w_3136_);
or (w_1322_, w_0240_, w_0967_);
and (w_0528_, w_0580_, w_1671_);
not (w_2269_, w_0911_);
or (w_2228_, w_1437_, w_1948_);
and (w_0898_, w_2959_, w_0407_);
not (w_0444_, w_2981_);
and (w_2638_, w_1844_, w_0439_);
or (w_0721_, w_1856_, w_2480_);
not (w_2921_, w_2808_);
or (w_1382_, w_1756_, w_3082_);
and (w_2651_, w_2236_, w_3212_);
and (w_0824_, in8[2], w_1533_);
and (out15[2], w_3410_, w_2643_);
and (w_1935_, w_0681_, w_0569_);
and (w_2861_, w_0004_, w_0166_);
and (w_2640_, w_0781_, w_1683_);
and (w_3511_, in9[6], in10[2]);
or (w_2027_, w_0688_, w_1300_);
not (w_0617_, in7[2]);
and (w_0037_, w_1345_, w_1430_);
or (w_0547_, w_2659_, w_0820_);
and (w_3420_, w_2806_, w_2143_);
not (w_0766_, w_0167_);
or (w_1522_, w_2560_, w_1049_);
and (w_3336_, in7[0], w_2023_);
and (w_2979_, w_2801_, w_0572_);
or (w_2983_, w_2450_, w_0515_);
and (w_0689_, w_0149_, w_1416_);
not (w_3000_, w_1248_);
not (w_1116_, w_2106_);
and (w_1166_, w_2935_, w_0338_);
and (w_1911_, w_3124_, w_1969_);
or (w_1823_, w_2552_, w_3146_);
and (w_1272_, w_2570_, w_3494_);
not (w_0145_, w_1867_);
and (w_3382_, w_1067_, w_0172_);
not (w_1434_, w_1026_);
and (w_2883_, w_2423_, w_1011_);
and (w_1586_, w_1535_, w_0271_);
and (w_2663_, w_1590_, w_2318_);
and (w_0216_, w_0265_, w_1951_);
and (w_1113_, w_0887_, w_0594_);
or (w_2427_, w_0374_, w_2919_);
and (w_2152_, w_2645_, w_1132_);
and (w_2326_, w_2959_, w_0671_);
or (w_2214_, w_0527_, w_3251_);
and (w_3510_, w_2739_, w_1109_);
or (w_0232_, w_1174_, w_0064_);
or (w_0098_, w_1105_, w_2116_);
or (w_1093_, w_3124_, w_0482_);
and (w_0473_, w_1275_, w_3292_);
not (w_0342_, w_0190_);
or (w_2138_, w_0349_, w_1692_);
and (w_0866_, in8[1], w_0552_);
and (w_2387_, w_0619_, w_1710_);
not (w_1486_, w_0220_);
or (w_1765_, w_0188_, w_1563_);
or (w_0928_, w_3352_, w_0271_);
not (w_0189_, w_1671_);
or (w_3183_, w_0596_, w_2191_);
and (w_0693_, w_2360_, w_2215_);
and (w_2066_, w_3385_, w_3039_);
or (out18[5], w_1969_, w_3330_);
and (w_2976_, w_2383_, w_3181_);
and (w_3309_, w_1474_, w_3175_);
not (w_0355_, w_1939_);
and (w_0235_, w_3405_, w_1535_);
or (w_1370_, w_3443_, w_3404_);
or (w_2772_, w_1069_, w_2846_);
not (w_0969_, w_2612_);
or (w_2178_, w_2935_, w_0338_);
and (w_0105_, in14[3], w_2744_);
not (w_0285_, w_0055_);
or (w_2615_, w_1888_, w_0854_);
and (w_1455_, w_1632_, w_1294_);
and (w_2844_, in14[3], in13[3]);
or (w_0746_, out14[0], out15[0]);
or (w_2776_, w_3412_, w_0804_);
and (w_0788_, w_0442_, w_2341_);
and (w_3438_, w_2153_, w_1323_);
not (w_0348_, w_2771_);
and (w_2313_, w_0728_, w_3311_);
and (w_1194_, w_2185_, w_1030_);
or (w_1928_, in15[0], w_0509_);
not (w_0479_, w_2417_);
and (w_1505_, w_0421_, w_1895_);
or (w_0449_, w_1926_, w_1446_);
and (w_1241_, w_1758_, w_1874_);
and (w_0129_, w_2125_, w_2232_);
or (w_3298_, w_1122_, w_1839_);
or (w_3506_, w_0436_, w_1448_);
and (w_3484_, in13[6], w_2556_);
or (w_1946_, in11[5], w_1984_);
and (w_0403_, w_2064_, w_3269_);
and (w_2417_, w_0380_, w_3524_);
and (w_1223_, w_0859_, w_1529_);
and (w_3423_, w_2196_, w_1641_);
or (w_0673_, w_3470_, w_2372_);
and (w_2970_, w_0857_, w_1512_);
not (w_3206_, w_2968_);
and (w_0872_, w_1567_, w_2080_);
not (w_1701_, w_0156_);
or (w_0979_, w_0249_, w_1643_);
or (w_2631_, w_3286_, w_0932_);
or (w_2477_, w_3308_, w_0467_);
or (w_3094_, w_0299_, w_3078_);
not (w_0365_, in4[4]);
not (w_2871_, w_0549_);
and (w_3194_, in13[1], w_2127_);
not (w_2194_, in3[1]);
not (w_2724_, w_1827_);
or (w_1608_, w_1435_, w_3133_);
or (w_2284_, w_0927_, w_1425_);
not (w_0538_, w_1963_);
and (w_3318_, w_2505_, w_0900_);
or (w_2359_, w_0839_, w_2432_);
not (w_1340_, w_2738_);
and (w_0978_, w_2873_, w_0717_);
and (w_0646_, w_3231_, w_0129_);
or (w_0028_, w_2028_, w_1426_);
and (w_2127_, w_2836_, w_1933_);
not (w_2592_, w_2728_);
and (w_2945_, w_0377_, w_1172_);
or (w_2354_, w_0666_, w_0271_);
not (w_0583_, w_1030_);
or (w_1813_, w_2137_, w_0174_);
not (w_1410_, w_1007_);
or (w_1943_, w_2098_, w_2875_);
or (w_0825_, w_0866_, w_2889_);
or (w_0908_, w_1753_, w_0523_);
not (w_3512_, w_1951_);
or (w_0109_, w_1629_, w_1441_);
and (out1[3], w_2706_, w_2805_);
or (w_2128_, w_3456_, w_3135_);
not (w_0840_, in4[3]);
and (w_0185_, w_2723_, w_0823_);
or (w_1230_, w_1660_, w_1347_);
and (w_3386_, w_3148_, w_1896_);
and (w_3221_, w_2353_, w_2109_);
and (w_0262_, w_1044_, w_2522_);
and (w_1183_, w_0277_, w_1085_);
and (w_0822_, w_2207_, w_2674_);
or (w_3397_, w_3445_, w_0650_);
and (w_0045_, w_1423_, w_0684_);
or (w_0618_, w_2283_, w_1592_);
and (w_0874_, w_0696_, w_2962_);
or (w_0602_, w_2578_, w_0155_);
not (w_0413_, w_2646_);
or (w_1524_, w_0895_, w_0460_);
not (w_2685_, in5[0]);
or (w_3299_, w_2712_, w_0919_);
not (w_1246_, w_1474_);
not (w_3137_, w_2503_);
and (w_0834_, w_0707_, w_0597_);
or (w_2823_, w_0864_, w_1288_);
or (w_1609_, w_2652_, w_0092_);
and (w_3479_, w_2937_, w_2953_);
and (w_1779_, w_1548_, w_1520_);
and (out2[4], w_2823_, w_2872_);
and (w_2421_, in15[4], w_3026_);
or (w_3067_, w_1436_, w_3040_);
or (w_2454_, w_1473_, w_2376_);
or (w_3211_, w_2105_, w_3369_);
not (w_1456_, w_3399_);
or (w_1672_, w_2128_, w_2956_);
and (w_0818_, w_2380_, w_0752_);
and (w_2732_, w_2455_, w_0031_);
and (w_0433_, w_1501_, w_1706_);
or (w_1038_, w_0049_, w_0121_);
and (w_0906_, w_1882_, w_1451_);
or (w_0172_, w_1290_, w_0876_);
or (w_1318_, w_3015_, w_1514_);
and (w_2978_, w_0117_, w_1693_);
or (w_0384_, in3[0], w_2940_);
or (w_2891_, w_1582_, w_1561_);
or (w_2649_, out13[6], w_3418_);
or (w_0981_, w_1407_, w_0344_);
and (w_3066_, in12[2], w_1461_);
not (w_0006_, w_1915_);
or (w_0195_, w_2563_, w_1399_);
or (w_0806_, w_2177_, w_2106_);
not (w_0909_, in6[2]);
or (out11[0], w_1151_, w_2378_);
and (w_1462_, w_2257_, w_0198_);
and (w_2832_, w_0781_, w_3348_);
and (w_0907_, out15[0], w_2803_);
not (w_1662_, w_0310_);
and (w_3038_, w_2868_, w_1525_);
and (w_1668_, w_0237_, w_2139_);
or (w_1866_, w_0192_, w_3125_);
or (w_3250_, w_2477_, w_3450_);
not (w_1428_, w_2642_);
and (w_3226_, w_0538_, w_1615_);
or (out19[3], w_0501_, w_1506_);
and (w_3402_, w_1027_, w_0779_);
not (w_1443_, in16[5]);
or (w_2484_, in6[2], in5[1]);
and (w_3287_, w_1339_, w_2218_);
and (w_1393_, w_0827_, w_0811_);
and (w_2504_, w_2601_, w_1906_);
and (w_1681_, w_3328_, w_0295_);
or (w_1089_, w_0970_, w_2112_);
or (w_2647_, w_1967_, w_2769_);
or (w_0719_, w_0463_, w_1124_);
or (w_0212_, w_1877_, w_0372_);
and (w_3178_, w_1368_, w_1955_);
or (w_2253_, w_2571_, w_0110_);
or (w_1726_, w_2564_, w_3130_);
not (w_0744_, w_2546_);
or (w_0976_, w_3007_, w_0834_);
or (w_2212_, w_3510_, w_1519_);
not (w_0019_, w_2601_);
and (w_0353_, w_3472_, w_1411_);
or (w_3356_, w_0989_, w_0033_);
and (w_1263_, w_0396_, w_2539_);
or (w_0691_, w_0034_, w_1621_);
or (w_2927_, w_1622_, w_2789_);
not (w_3345_, in15[0]);
or (w_3025_, w_3498_, w_3518_);
or (w_1502_, in7[3], w_1745_);
and (w_1499_, w_3154_, w_3467_);
and (w_2118_, w_1529_, w_1908_);
and (w_0833_, w_0289_, w_2272_);
and (out14[4], w_2779_, w_2866_);
not (w_3327_, w_0344_);
and (w_2894_, w_0808_, w_1920_);
or (w_0248_, w_0609_, w_2468_);
and (w_2518_, w_2237_, w_2756_);
not (w_0764_, w_0867_);
or (w_1956_, w_3328_, w_0295_);
and (w_2292_, w_3002_, w_0503_);
not (w_0222_, w_1191_);
and (w_0057_, w_2371_, w_1320_);
or (w_2275_, w_0720_, w_2490_);
not (w_1557_, w_3090_);
or (w_0916_, w_1981_, w_0715_);
or (w_0247_, w_2465_, w_2700_);
not (w_3491_, in6[1]);
or (w_0272_, w_0909_, w_0098_);
or (w_2462_, w_2153_, w_1323_);
not (w_0683_, w_3220_);
or (out5[5], w_1997_, w_2240_);
or (w_0315_, w_0831_, w_3202_);
and (w_3404_, w_1200_, w_1353_);
not (w_1452_, w_3021_);
not (w_1210_, in11[3]);
and (w_0465_, w_2073_, w_1495_);
or (w_0887_, w_2910_, w_3427_);
or (w_3150_, w_2761_, w_2597_);
or (w_0230_, w_0323_, w_1959_);
and (w_0300_, w_1007_, w_2230_);
and (w_0299_, w_1680_, w_1181_);
or (w_3131_, w_2175_, w_0693_);
or (out20[3], w_0227_, w_0367_);
not (w_2088_, w_1148_);
and (w_3093_, w_1419_, w_1993_);
or (w_0351_, w_0337_, w_2385_);
or (out18[0], w_0666_, w_3297_);
not (w_0772_, in5[5]);
or (w_0873_, w_0403_, w_1647_);
or (w_0361_, w_0446_, w_3204_);
not (w_2019_, w_2518_);
not (w_1402_, w_2907_);
and (w_3418_, w_1673_, w_1969_);
or (w_1910_, w_2198_, w_3206_);
and (w_0687_, in12[3], w_1748_);
or (w_1075_, w_2788_, w_2323_);
or (w_0531_, w_2281_, w_2718_);
and (w_0555_, in1[1], in2[1]);
or (w_2781_, w_1774_, w_2845_);
and (w_2246_, in14[2], in13[2]);
and (w_2788_, w_0550_, w_1150_);
or (w_0254_, w_1753_, w_2602_);
or (w_1128_, w_1314_, w_0554_);
or (w_0233_, w_2474_, w_0064_);
and (w_0967_, w_1877_, w_1761_);
not (w_2386_, w_1835_);
not (w_3128_, w_1263_);
or (w_0530_, w_1736_, w_0794_);
and (w_2703_, w_1202_, w_3145_);
not (w_2073_, w_1535_);
and (w_0469_, in3[2], w_3303_);
not (w_0724_, w_1406_);
or (w_2136_, w_3073_, w_3306_);
and (w_0659_, w_0599_, w_0489_);
and (w_0033_, w_2108_, w_2201_);
and (w_2497_, w_2936_, w_1367_);
and (w_0757_, w_3248_, w_2427_);
and (w_2627_, in7[1], w_3163_);
or (out8[4], w_3207_, w_0656_);
and (w_1962_, w_0734_, w_1379_);
and (w_0066_, w_0550_, w_3374_);
not (w_0380_, w_2028_);
or (w_2160_, w_0020_, w_0585_);
and (w_2085_, w_2310_, w_0867_);
and (w_0176_, w_0871_, w_1699_);
not (w_0929_, w_2132_);
and (w_1063_, w_2512_, w_1760_);
or (w_0281_, w_1330_, w_3198_);
not (w_0963_, in4[1]);
or (w_2220_, w_0370_, w_0577_);
or (w_2134_, w_0086_, w_3370_);
not (w_0850_, w_2484_);
and (w_0615_, in15[3], in16[3]);
not (w_1315_, in14[5]);
and (w_1478_, w_1015_, w_2981_);
or (w_1178_, w_0531_, w_2252_);
or (w_1090_, w_2819_, w_1052_);
and (w_0817_, w_3096_, w_0419_);
or (out19[4], w_2474_, w_1232_);
or (w_1103_, out9[0], w_2968_);
and (w_1483_, w_3019_, w_1068_);
or (w_1389_, in6[5], w_1664_);
and (w_2666_, w_1372_, w_0184_);
or (w_0441_, w_0601_, w_1404_);
and (w_2040_, w_3474_, w_1185_);
not (w_1317_, in12[0]);
or (w_2035_, w_0873_, w_1022_);
and (w_0168_, w_2356_, w_1047_);
and (w_0591_, w_0551_, w_2488_);
or (w_1824_, w_2910_, w_2596_);
or (w_3027_, in3[2], w_3280_);
or (w_0716_, in15[7], w_2764_);
not (w_3378_, w_1907_);
and (w_1790_, w_1418_, w_1568_);
or (w_2250_, w_0708_, w_2947_);
or (w_0725_, w_1699_, w_0455_);
and (w_0147_, w_3424_, w_1645_);
not (w_3362_, w_2556_);
not (w_0515_, w_1454_);
or (w_1854_, w_0943_, w_2656_);
and (w_2216_, w_3387_, w_1672_);
or (w_0653_, w_2411_, w_2815_);
or (w_2783_, w_0370_, w_1239_);
not (w_3151_, in16[6]);
not (w_3374_, w_3430_);
and (w_2958_, w_2314_, w_3077_);
and (w_1066_, w_2175_, w_0418_);
and (w_1088_, w_2931_, w_2810_);
or (w_0588_, w_1026_, w_1267_);
and (w_2558_, w_0427_, w_2664_);
not (w_0368_, w_3119_);
and (w_1537_, w_1676_, w_2739_);
and (w_1748_, w_1542_, w_1167_);
and (w_3168_, w_1519_, w_2057_);
and (w_2768_, w_1463_, w_2767_);
and (w_0856_, w_2451_, w_0899_);
and (w_0821_, w_2506_, w_1074_);
not (w_3515_, w_2568_);
or (w_2112_, w_0024_, w_0732_);
or (w_2734_, in4[1], w_2327_);
and (w_1963_, w_1892_, w_3314_);
and (w_1239_, w_0215_, w_2434_);
or (w_0047_, w_2049_, w_0190_);
or (w_0162_, w_1354_, w_1070_);
and (w_3059_, w_2631_, w_3419_);
not (w_0042_, w_1118_);
and (w_3422_, w_1093_, w_3235_);
or (w_0224_, w_0102_, w_1467_);
not (w_1404_, out13[0]);
and (w_1016_, w_2508_, w_1318_);
and (w_2364_, in9[6], in10[6]);
or (w_0728_, w_1210_, w_0813_);
and (w_0858_, w_0240_, w_2324_);
or (w_2041_, in13[4], w_0259_);
and (w_2345_, w_0063_, w_3387_);
not (w_2469_, w_1689_);
and (out21[2], w_2522_, w_0886_);
or (w_1567_, w_3139_, w_1985_);
or (w_0512_, w_3005_, w_0914_);
not (w_1313_, w_0774_);
and (w_1633_, w_0329_, w_0154_);
not (w_1302_, w_1310_);
and (w_0567_, w_0543_, w_0230_);
or (w_2272_, w_1878_, w_2274_);
and (w_1533_, w_0795_, w_2890_);
not (w_3236_, w_2244_);
or (w_1958_, w_3316_, w_0330_);
and (w_1138_, w_3220_, w_0744_);
not (w_0081_, w_0743_);
and (w_3333_, in7[3], w_1745_);
and (w_1095_, w_0207_, w_0058_);
not (w_1039_, w_3230_);
and (w_1108_, in13[4], w_0259_);
or (w_2501_, w_2646_, w_3413_);
not (w_0667_, w_0877_);
and (w_0275_, in4[4], w_1611_);
or (w_2723_, w_2882_, w_1099_);
or (w_1165_, w_1211_, w_2633_);
or (w_3109_, w_3442_, w_1952_);
and (w_1207_, w_0035_, w_1269_);
and (w_1599_, w_2858_, w_2313_);
or (w_2540_, w_0007_, w_2525_);
and (w_3132_, w_0358_, w_3008_);
and (w_3050_, w_1665_, w_1129_);
or (w_2080_, w_0010_, w_3392_);
or (w_0016_, w_1365_, w_3166_);
and (w_0507_, w_0225_, w_1333_);
not (w_0527_, w_1843_);
and (w_0086_, w_1494_, w_2776_);
or (w_2308_, w_2304_, w_0468_);
not (w_3437_, w_1944_);
and (w_1922_, w_0682_, w_1125_);
and (w_2932_, w_2533_, w_1478_);
and (w_1203_, w_0148_, w_3528_);
not (w_1249_, w_3321_);
and (w_1648_, in15[1], w_1213_);
or (w_2144_, w_0337_, w_2668_);
not (w_0359_, w_1780_);
and (out2[0], w_0962_, w_1021_);
or (w_2729_, w_2358_, w_0695_);
and (w_0404_, w_0036_, w_0855_);
or (w_0684_, w_2086_, w_3528_);
or (w_3008_, w_1835_, w_1439_);
or (w_2813_, in1[0], in2[1]);
and (w_3214_, w_1628_, w_2396_);
and (w_0426_, w_2708_, w_0930_);
or (w_1578_, w_0646_, w_2816_);
and (w_0810_, w_1931_, w_0078_);
or (w_3315_, w_2958_, w_0938_);
or (w_2645_, w_1361_, w_1187_);
or (w_2368_, w_0372_, w_2270_);
and (w_0214_, w_0944_, w_0787_);
and (w_2487_, w_2935_, w_0873_);
and (out2[2], w_2983_, w_1341_);
and (w_0711_, w_2444_, w_2860_);
not (w_0753_, w_0779_);
or (w_0018_, w_1948_, w_2894_);
or (w_2132_, w_2167_, w_2344_);
and (w_1005_, w_1835_, w_1439_);
not (w_2107_, in13[5]);
or (w_3387_, w_2531_, w_1075_);
or (w_2966_, w_2716_, w_1453_);
or (w_3114_, w_3040_, w_1401_);
or (w_0902_, w_1947_, w_0660_);
and (w_2571_, w_1291_, w_1322_);
not (w_1558_, w_2422_);
or (w_1827_, in6[1], in5[0]);
or (w_3354_, w_3396_, w_0250_);
and (w_2281_, in5[1], w_0692_);
and (w_3324_, w_3248_, w_0755_);
and (w_3202_, w_0000_, w_3107_);
or (w_3144_, in1[1], in2[1]);
or (out1[5], w_1772_, w_3418_);
or (w_2347_, w_3058_, w_1148_);
and (w_0540_, w_0826_, w_0741_);
and (w_0487_, w_0322_, w_2371_);
and (out7[2], w_2695_, w_2138_);
or (w_1292_, w_0956_, w_0385_);
or (w_1474_, w_2758_, w_0750_);
or (w_0132_, w_1900_, w_2492_);
and (w_2369_, in6[3], in5[2]);
not (w_0107_, w_0629_);
or (w_3433_, w_0275_, w_1447_);
and (out17[6], w_1429_, w_1714_);
and (w_1771_, w_0742_, w_2253_);
or (w_3452_, w_0971_, w_1215_);
not (w_1879_, w_3429_);
or (w_3441_, w_0106_, w_1497_);
or (w_1568_, w_2263_, w_2909_);
or (w_3165_, w_3247_, w_3227_);
and (w_2771_, w_2078_, w_3131_);
or (w_1438_, w_2787_, w_3346_);
or (w_1774_, w_0952_, w_2896_);
or (w_0780_, w_3494_, w_0935_);
or (w_2905_, w_1207_, w_2264_);
or (w_2455_, w_3073_, w_1023_);
and (out21[0], w_0113_, w_2530_);
and (w_1197_, w_3444_, w_3366_);
not (w_2021_, w_0159_);
and (w_2989_, w_2173_, w_3068_);
and (w_3060_, w_2905_, w_0620_);
and (w_2847_, w_0988_, w_1803_);
and (w_3091_, w_1217_, w_3080_);
or (w_2586_, w_2932_, w_2989_);
or (w_0849_, w_3267_, w_2820_);
and (w_0762_, w_1504_, w_1736_);
or (w_2779_, w_3285_, w_0570_);
not (w_2046_, in9[1]);
or (w_0501_, w_0347_, w_1863_);
and (w_0446_, w_0322_, w_2778_);
or (w_3317_, w_2563_, w_1616_);
and (w_2340_, w_3294_, w_2592_);
or (w_1036_, w_3081_, w_0432_);
and (w_2856_, w_2292_, w_2979_);
or (w_1639_, w_3191_, w_2110_);
not (w_0570_, w_2004_);
not (w_0931_, w_2626_);
and (w_1811_, w_0305_, w_1975_);
and (w_2662_, w_1095_, w_2073_);
and (w_1953_, w_2432_, w_3142_);
and (w_0533_, w_0310_, w_0320_);
and (w_1643_, w_3494_, w_2959_);
not (w_2689_, w_0378_);
or (w_1264_, w_3473_, w_1833_);
or (w_0063_, w_1442_, w_1466_);
or (w_1459_, w_3048_, w_2102_);
not (w_2807_, w_1365_);
and (w_2478_, w_0133_, w_1832_);
not (w_1805_, in14[3]);
and (w_0666_, w_0705_, w_1405_);
and (w_1035_, out14[0], out15[0]);
or (w_2825_, w_2959_, w_2667_);
or (w_1372_, w_0452_, w_1516_);
or (w_2784_, w_2935_, w_3051_);
or (w_2115_, w_1317_, w_2675_);
or (w_3507_, w_2703_, w_2154_);
not (w_3316_, in12[1]);
and (out17[3], w_0804_, w_3021_);
or (w_1071_, w_2879_, w_1480_);
and (w_0604_, w_1007_, w_0411_);
and (w_2460_, in15[6], in16[6]);
and (w_0656_, w_2959_, w_0217_);
or (w_1579_, out14[4], w_2923_);
or (w_1193_, w_0035_, w_2356_);
or (w_2304_, w_2515_, w_2755_);
and (w_1604_, w_1725_, w_0686_);
and (w_0414_, w_0994_, w_3244_);
and (w_1678_, w_2565_, w_0431_);
not (w_3198_, w_0939_);
or (w_2597_, w_0301_, w_1309_);
not (w_2312_, w_2435_);
and (w_2881_, in11[1], w_0965_);
and (w_2036_, w_0217_, w_1080_);
and (out22[1], w_3428_, w_3239_);
and (w_0337_, in5[3], w_3460_);
or (w_2774_, w_0469_, w_0576_);
or (w_0645_, w_2064_, w_2504_);
or (out12[4], w_1270_, w_2203_);
or (w_0135_, w_0840_, w_2441_);
and (w_2309_, w_2772_, w_0267_);
or (out20[2], w_1400_, w_2960_);
and (w_1686_, w_3037_, w_0298_);
not (w_2439_, w_2940_);
or (w_1037_, w_0217_, w_0244_);
not (w_1695_, w_3384_);
and (w_1845_, w_0034_, w_2073_);
or (w_2740_, w_1479_, w_0219_);
and (w_2843_, w_0572_, w_2749_);
or (out3[2], w_1391_, w_1177_);
or (w_2920_, w_0545_, w_1191_);
and (w_0015_, w_0802_, w_3297_);
or (w_1882_, w_3367_, w_0245_);
or (w_3467_, w_2851_, w_2939_);
or (w_2475_, in3[1], w_0830_);
and (w_3193_, w_1436_, w_3497_);
and (w_0372_, w_1776_, w_0366_);
or (w_0274_, w_1250_, w_2251_);
and (w_3181_, w_1456_, w_1583_);
and (w_1332_, w_0128_, w_0412_);
or (w_1248_, in13[3], w_3323_);
or (w_2748_, w_2316_, w_0293_);
or (w_2812_, in3[4], w_2699_);
or (w_0294_, w_0105_, w_3515_);
and (w_3466_, w_1918_, w_2585_);
or (w_3454_, w_2393_, w_1629_);
and (w_2678_, w_3310_, w_2624_);
not (w_1580_, w_2361_);
and (w_0078_, w_0673_, w_0218_);
or (w_1602_, w_1747_, w_1095_);
or (w_2011_, in9[7], in10[7]);
or (w_0921_, w_0506_, w_1472_);
or (w_1545_, w_2185_, w_0669_);
or (w_0614_, w_3377_, w_3049_);
or (w_2866_, w_2991_, w_2004_);
not (w_1433_, w_2992_);
not (w_3140_, w_1507_);
not (w_3501_, w_1174_);
and (w_1885_, w_2712_, w_1728_);
or (w_1778_, w_1616_, w_3174_);
and (w_3297_, w_3063_, w_2757_);
or (w_2681_, w_0034_, w_0322_);
and (w_3369_, w_2652_, w_0092_);
not (w_1860_, w_1097_);
or (w_1680_, w_2283_, w_1326_);
or (w_3448_, w_2101_, w_0890_);
or (w_1112_, w_1849_, out16[7]);
not (w_1529_, w_2961_);
or (w_2929_, w_1843_, w_2623_);
or (w_3370_, w_1515_, w_1585_);
and (w_0685_, in7[2], w_1311_);
or (w_1788_, w_0694_, w_0170_);
or (w_0400_, in8[2], w_1851_);
and (w_2146_, w_0966_, w_2147_);
and (w_3061_, w_3033_, w_1445_);
not (w_2560_, in6[4]);
or (w_1925_, w_0139_, w_2489_);
not (w_1024_, in15[6]);
not (w_1969_, w_3352_);
not (w_0104_, in12[4]);
and (w_3127_, w_0438_, w_1163_);
or (w_0251_, w_2924_, w_2564_);
and (w_0322_, w_2962_, w_2503_);
and (w_2576_, w_0580_, w_0457_);
not (w_2702_, w_0297_);
and (w_2537_, w_1788_, w_2762_);
and (w_0786_, w_0322_, w_2153_);
and (w_2719_, w_0722_, w_3270_);
and (w_2950_, w_1674_, w_0528_);
or (w_2335_, w_0055_, w_1305_);
and (w_0171_, w_0729_, w_1268_);
and (w_2629_, w_1806_, w_0261_);
not (w_0174_, w_0196_);
and (w_0059_, w_1616_, w_3174_);
or (w_0071_, w_1737_, w_3105_);
or (w_0116_, w_2394_, w_2536_);
not (w_1786_, w_2313_);
not (w_1466_, w_1150_);
or (w_0752_, w_0383_, w_0150_);
not (w_0273_, w_0232_);
and (out13[3], w_2706_, w_2805_);
and (w_0205_, w_0849_, w_0386_);
and (w_1391_, w_1150_, w_1380_);
or (w_3023_, w_0178_, w_1599_);
not (w_3367_, in11[5]);
not (w_0100_, w_3187_);
or (w_2446_, w_1477_, w_0513_);
not (w_1636_, w_1479_);
or (w_0642_, w_3152_, w_0085_);
and (w_1242_, w_0928_, w_1006_);
or (out24[0], w_1035_, w_2775_);
or (w_1952_, w_0582_, w_0325_);
or (w_0982_, w_1149_, w_0236_);
and (w_2452_, in12[1], w_2943_);
or (w_2674_, w_0758_, w_0578_);
or (w_0263_, w_1949_, w_2820_);
not (w_0227_, w_1188_);
or (w_1509_, w_0659_, w_3463_);
or (w_2643_, w_3328_, w_1304_);
and (w_1495_, w_0493_, w_2337_);
and (w_3012_, w_1986_, w_0195_);
and (w_1873_, w_2484_, w_2300_);
and (w_0851_, w_3397_, w_3219_);
or (w_1785_, w_3477_, w_2999_);
and (w_1419_, in1[0], in2[0]);
not (w_1430_, w_0663_);
or (w_1598_, w_3194_, w_0559_);
not (w_2291_, w_2840_);
not (w_3520_, w_2542_);
and (w_1732_, w_3100_, w_0885_);
and (w_2680_, w_2560_, w_1049_);
and (w_0269_, w_2645_, w_3507_);
and (w_3171_, w_3339_, w_2874_);
and (w_0599_, w_0725_, w_1649_);
or (w_3389_, w_2494_, w_1899_);
not (w_1705_, w_0510_);
or (w_0697_, w_0365_, w_1886_);
and (w_1439_, w_0961_, w_1293_);
or (out8[2], w_1620_, w_0015_);
and (w_3158_, w_0738_, w_0981_);
not (w_0329_, in4[5]);
not (w_0595_, w_2899_);
or (w_0239_, w_2858_, w_2313_);
and (w_1475_, w_2086_, w_2827_);
and (w_2468_, w_2073_, w_3292_);
and (w_1460_, w_0793_, w_0279_);
and (w_1841_, w_0020_, w_0585_);
or (w_0466_, w_1735_, w_0153_);
and (w_0876_, w_3405_, w_2570_);
or (out20[4], w_2120_, w_0283_);
or (w_1176_, w_3288_, w_1762_);
and (w_1610_, w_0217_, w_0336_);
or (out5[2], w_1845_, w_2599_);
and (out16[0], w_0633_, w_2664_);
and (w_2480_, w_1593_, w_1031_);
and (w_2188_, w_1038_, w_1193_);
and (w_2799_, w_1146_, w_3305_);
and (w_2224_, w_3242_, w_0838_);
or (w_0334_, in16[6], w_2907_);
not (w_0771_, w_1230_);
or (w_1780_, in11[2], w_1703_);
and (w_3268_, w_3492_, w_2526_);
not (w_1335_, w_3323_);
not (w_0805_, w_2695_);
and (w_0288_, w_1942_, w_0345_);
and (w_1034_, out14[5], w_1761_);
and (w_0524_, w_2093_, w_3032_);
and (w_2222_, w_1442_, w_3430_);
or (w_2002_, w_2995_, w_2331_);
or (w_0108_, w_0622_, w_1633_);
or (w_2984_, w_3465_, w_3161_);
not (w_3264_, in7[0]);
or (w_1590_, w_0617_, w_1055_);
and (w_1647_, w_1853_, w_1791_);
or (w_2287_, w_1263_, w_2611_);
and (out6[2], w_1474_, w_1141_);
or (w_0857_, in1[4], in2[5]);
and (w_0253_, w_1393_, w_0056_);
and (w_1277_, w_0562_, w_1976_);
or (w_2860_, w_2726_, w_1988_);
or (w_1973_, w_3112_, w_0262_);
or (w_2184_, w_1016_, w_2219_);
or (w_0671_, w_0680_, w_1087_);
or (w_1394_, w_3527_, w_2150_);
or (w_1060_, in15[5], w_2100_);
and (out24[2], w_1929_, w_0920_);
and (w_3291_, w_0379_, w_0029_);
and (w_0623_, w_2365_, w_3462_);
and (w_2878_, w_2512_, w_0445_);
and (w_1399_, w_2334_, w_3347_);
and (w_3233_, w_2765_, w_2521_);
or (w_0705_, w_1747_, w_0464_);
and (w_0971_, in8[3], w_1397_);
and (w_1942_, w_3436_, w_1996_);
or (w_0966_, w_3491_, w_0702_);
and (w_0539_, w_1853_, w_1969_);
not (w_0964_, w_3059_);
and (w_2262_, w_0553_, w_1918_);
not (w_2614_, w_3297_);
or (w_0154_, w_0577_, w_0397_);
not (w_1384_, w_1399_);
and (w_2431_, w_1134_, w_0756_);
or (w_1844_, w_0105_, w_0621_);
not (w_3364_, w_1344_);
or (w_0186_, w_0214_, w_2803_);
or (w_0161_, w_2982_, w_0901_);
or (w_1070_, w_2665_, w_0026_);
or (w_1157_, w_1498_, w_3075_);
and (w_1795_, w_1942_, out16[3]);
and (w_0518_, w_2005_, w_3136_);
and (w_2542_, in1[3], in2[4]);
not (w_1386_, w_2619_);
and (w_3218_, w_1656_, w_0224_);
and (w_1503_, w_3021_, w_0482_);
not (w_0638_, w_1766_);
or (w_1168_, w_1410_, w_0602_);
or (w_3355_, w_0240_, w_2324_);
or (w_1163_, w_3505_, w_1421_);
or (w_1083_, w_1482_, w_2330_);
not (w_1682_, w_1976_);
or (w_1114_, w_1605_, w_2577_);
and (w_2531_, w_2461_, w_1723_);
and (w_2808_, w_3213_, w_1184_);
or (w_2790_, w_1320_, w_3337_);
not (w_0242_, w_0509_);
or (w_0790_, w_1743_, w_3224_);
and (w_0853_, w_2609_, w_0319_);
not (w_0532_, w_2844_);
or (w_1847_, w_2449_, w_3095_);
not (w_0415_, w_1679_);
and (w_2547_, w_2935_, w_2180_);
not (w_1218_, w_1471_);
not (w_3161_, w_0425_);
or (w_1689_, w_2935_, w_2180_);
and (w_1650_, w_1740_, w_0635_);
or (w_0735_, w_0269_, w_3402_);
not (w_0815_, w_0311_);
not (w_1710_, w_1342_);
or (w_3217_, w_3452_, w_1912_);
not (w_1366_, in6[3]);
and (w_3292_, w_1602_, w_1545_);
or (w_0362_, w_1967_, w_1328_);
and (out21[5], w_2341_, w_2259_);
or (w_1009_, in15[3], w_1618_);
or (w_3527_, w_1555_, w_3022_);
or (w_3283_, w_1654_, w_2848_);
or (w_2237_, w_2926_, w_3064_);
and (w_1592_, w_0099_, w_1449_);
or (w_2330_, w_2982_, w_1221_);
and (w_2393_, w_0034_, w_2961_);
or (w_0813_, w_1573_, w_0300_);
and (w_3015_, w_1434_, w_3357_);
or (w_0801_, w_1844_, w_0439_);
or (w_2930_, w_3034_, w_1737_);
or (w_2736_, w_1927_, w_1783_);
and (w_2067_, w_3149_, w_2220_);
or (w_3262_, w_0889_, w_2076_);
or (w_2942_, w_2413_, w_0736_);
or (w_2257_, w_2780_, w_2117_);
or (w_0613_, w_0496_, w_0014_);
and (w_2802_, w_1016_, w_2219_);
and (w_3130_, w_2465_, w_2700_);
or (w_1320_, w_1457_, w_2818_);
or (w_1857_, w_0501_, w_0173_);
not (w_1472_, w_0409_);
or (w_3020_, w_3154_, w_3467_);
or (out5[1], w_1911_, w_1887_);
or (w_2464_, w_0284_, w_2426_);
or (w_0418_, w_2174_, w_2710_);
and (w_1670_, w_2371_, w_1791_);
and (w_1003_, w_0894_, w_1711_);
not (w_2323_, w_1782_);
not (w_2985_, w_1504_);
not (w_1638_, w_0564_);
and (w_0985_, w_0778_, w_2025_);
or (w_2899_, w_1737_, w_0237_);
and (w_1891_, w_0048_, w_1261_);
or (w_2260_, w_2668_, w_2534_);
not (w_0759_, w_2536_);
or (w_0791_, w_0223_, w_2987_);
or (w_1287_, w_2156_, w_0743_);
and (w_0901_, w_0522_, w_1831_);
not (w_1396_, w_1754_);
or (w_3244_, w_3492_, w_2961_);
and (w_1262_, w_2416_, w_0228_);
and (w_0760_, w_1541_, w_2743_);
or (w_2803_, w_3031_, w_2315_);
or (w_1745_, w_1422_, w_1244_);
or (w_0991_, w_0416_, w_3292_);
and (w_2602_, w_1383_, w_0274_);
or (w_2805_, w_0804_, w_3510_);
and (out17[1], w_1737_, w_0658_);
and (w_0183_, w_1141_, w_3492_);
and (w_2016_, w_1605_, w_3089_);
or (w_1593_, w_3085_, w_1994_);
and (w_3329_, w_0584_, w_2338_);
and (out4[2], w_3055_, w_0806_);
or (w_3276_, in14[6], w_3103_);
and (w_0393_, w_0772_, w_1189_);
and (w_3509_, w_0873_, w_1022_);
and (w_1450_, w_0666_, w_2343_);
not (w_1655_, out15[0]);
and (w_1903_, w_2086_, w_3218_);
and (w_1775_, w_1366_, w_2260_);
and (w_1874_, w_1114_, w_1298_);
and (w_0870_, in16[6], w_2907_);
or (w_1467_, w_1048_, w_0070_);
not (w_1863_, w_0723_);
or (w_0859_, w_0126_, w_2948_);
or (w_0143_, w_3438_, w_0199_);
not (w_1923_, w_2609_);
and (w_2357_, w_0586_, w_1009_);
and (w_3069_, w_2149_, w_0537_);
and (w_1283_, w_2009_, w_2266_);
and (w_3223_, w_0840_, w_2441_);
or (w_2334_, w_1858_, w_1712_);
not (w_1501_, in5[1]);
and (w_1191_, w_2825_, w_2165_);
not (w_0560_, w_0287_);
and (w_0508_, w_0363_, w_2249_);
or (w_0668_, in7[0], w_3090_);
or (w_3180_, w_2247_, w_1960_);
and (w_2003_, w_0942_, w_3501_);
and (w_2884_, w_1673_, w_1174_);
or (w_1031_, in12[6], w_3061_);
or (w_2505_, w_2107_, w_1357_);
and (w_0370_, in3[5], w_2195_);
or (w_3278_, w_2918_, w_0323_);
not (w_2015_, w_2887_);
not (w_2820_, w_3183_);
or (w_0148_, w_2800_, w_2400_);
or (w_1666_, w_3205_, w_2741_);
or (w_2039_, w_2713_, w_1786_);
or (w_2773_, w_0477_, w_3362_);
and (w_1913_, w_0252_, out13[3]);
or (w_1304_, w_2210_, w_1433_);
and (w_1890_, in4[3], w_1205_);
not (w_2104_, w_1752_);
and (w_2716_, w_2136_, w_3044_);
not (w_0435_, w_2838_);
or (w_0905_, w_2848_, w_1739_);
and (w_1888_, w_2618_, w_1604_);
and (w_0421_, w_1955_, w_0164_);
and (w_0984_, w_0005_, w_0313_);
and (out1[2], w_2050_, w_3117_);
and (w_0115_, w_2343_, w_1769_);
not (w_0587_, w_3291_);
and (w_2741_, w_1856_, w_2480_);
or (w_2062_, w_1369_, w_2221_);
or (w_1057_, w_2729_, w_2453_);
not (w_1078_, w_1609_);
or (w_2133_, out14[1], w_3172_);
or (w_1368_, w_0550_, w_2381_);
and (w_2728_, w_2064_, w_3352_);
or (w_0313_, w_1141_, w_2171_);
and (w_2438_, w_1915_, w_2425_);
and (w_0675_, w_3139_, w_1985_);
and (w_1100_, out14[1], w_3172_);
and (w_1244_, in6[4], in5[3]);
or (w_1496_, w_1463_, w_0234_);
or (w_1996_, w_0599_, w_1519_);
not (w_0802_, w_1393_);
not (w_1572_, w_3420_);
or (w_3270_, w_1773_, w_3519_);
and (w_1560_, w_0726_, w_3035_);
and (w_2306_, w_1455_, w_2543_);
and (w_2476_, w_1932_, w_3053_);
not (w_2766_, w_2011_);
or (w_3019_, w_1805_, w_1603_);
or (w_2337_, w_0550_, w_0999_);
not (w_1587_, w_3171_);
or (w_0013_, w_0000_, w_3107_);
and (w_2609_, w_3034_, w_3528_);
not (w_0079_, w_0390_);
and (w_3459_, w_0202_, w_0679_);
and (w_2151_, w_1698_, w_3321_);
or (w_0302_, w_2517_, w_0448_);
and (w_1862_, w_3165_, w_0353_);
not (w_2329_, w_3432_);
not (w_3421_, w_2656_);
or (w_1175_, w_1242_, w_0583_);
or (w_1278_, in9[7], in10[3]);
or (w_0025_, w_0421_, w_2338_);
or (w_1073_, w_3218_, w_2600_);
not (w_0679_, w_2369_);
or (w_0169_, w_2067_, w_0356_);
or (w_0231_, w_3358_, w_0832_);
or (w_2083_, w_2853_, w_1682_);
or (w_2055_, w_0322_, w_2371_);
or (w_1542_, w_2414_, w_1634_);
and (w_2254_, in7[2], w_2752_);
and (out6[0], w_3492_, w_0214_);
not (w_1027_, w_1746_);
and (w_0782_, w_2574_, w_1046_);
not (w_1387_, w_0250_);
or (w_1576_, w_1463_, out16[6]);
or (w_3351_, w_1888_, w_2867_);
and (w_2620_, w_0049_, w_0121_);
and (out22[2], w_0375_, w_0011_);
and (w_1573_, w_1410_, w_0602_);
and (w_3350_, w_0676_, w_1709_);
or (w_2467_, w_0346_, w_0797_);
or (w_0940_, w_2233_, w_2437_);
and (w_2191_, w_1560_, w_0583_);
or (w_0647_, w_1961_, w_2766_);
or (w_1782_, w_0550_, w_1150_);
or (w_2258_, in3[1], w_2666_);
or (w_0495_, w_0396_, w_2539_);
or (w_3481_, w_1259_, w_0486_);
and (w_0839_, w_2204_, w_2466_);
or (w_1186_, in16[7], w_1462_);
or (w_2491_, w_0479_, w_3304_);
and (w_1899_, w_0973_, w_2524_);
or (w_0823_, w_1337_, w_1219_);
and (w_0209_, w_1969_, w_0873_);
or (out12[2], w_2033_, w_2118_);
and (w_0237_, w_1904_, w_1319_);
and (w_3159_, out14[4], w_2923_);
not (w_2189_, w_3265_);
or (w_1625_, w_0343_, w_2016_);
and (w_2816_, w_2520_, w_1388_);
not (w_1994_, w_3061_);
not (w_1734_, out16[3]);
or (w_3234_, w_2194_, w_0194_);
or (w_1660_, w_3070_, w_2833_);
and (w_1664_, w_1212_, w_2797_);
not (w_2059_, in16[1]);
or (w_1219_, w_2514_, w_0869_);
not (w_2880_, w_3092_);
or (w_0166_, in5[5], w_0975_);
or (w_1153_, w_0800_, w_3351_);
and (w_1550_, w_1150_, w_2083_);
and (w_2362_, w_0943_, w_1519_);
or (out3[5], w_1897_, w_1759_);
not (w_2140_, w_2566_);
or (w_1225_, w_1552_, w_1158_);
and (w_0950_, w_1081_, w_1653_);
and (w_3013_, w_2078_, w_0629_);
not (w_2493_, w_2578_);
and (w_3243_, in4[1], w_1732_);
not (w_2661_, w_1770_);
or (w_2747_, w_2518_, w_1737_);
and (out4[4], w_0386_, w_1285_);
or (w_2605_, w_1876_, w_3183_);
not (w_2683_, w_0375_);
not (w_0718_, w_0321_);
and (w_2581_, w_2618_, w_2042_);
and (w_2798_, w_1286_, w_1799_);
or (w_1015_, w_2517_, w_3248_);
not (w_0889_, in3[2]);
or (w_3417_, w_1346_, w_2954_);
or (w_1029_, w_1095_, w_0408_);
and (w_0423_, w_3283_, w_2070_);
and (out15[1], w_2992_, w_2238_);
or (w_2836_, w_0082_, w_3312_);
and (w_2267_, w_2244_, w_0727_);
not (w_2617_, w_2481_);
and (w_0590_, in1[2], in2[3]);
and (w_1059_, w_0290_, w_2355_);
and (w_1446_, w_2677_, w_3221_);
or (w_2717_, w_2514_, w_3320_);
or (w_3057_, w_1359_, w_0784_);
or (w_0405_, w_0273_, w_2553_);
not (w_1924_, in16[3]);
or (out13[7], w_1279_, w_2092_);
and (w_0504_, w_3164_, w_3129_);
or (w_1274_, w_2832_, w_2040_);
not (w_2608_, w_0777_);
or (w_3474_, w_3197_, w_0107_);
not (w_0633_, w_0520_);
or (w_2568_, in14[3], w_2744_);
or (w_2296_, w_1466_, w_0583_);
or (w_2686_, w_3106_, w_3350_);
not (w_1773_, w_3469_);
and (w_3399_, w_1562_, w_0936_);
or (w_2280_, w_1474_, w_0271_);
or (w_2677_, w_2077_, w_2483_);
not (w_1548_, w_2067_);
or (w_0425_, in13[2], w_1807_);
or (w_2565_, w_2763_, w_0362_);
or (w_2076_, w_3210_, w_3514_);
not (w_3304_, w_3461_);
and (w_0835_, w_2518_, w_2667_);
and (w_3447_, w_2478_, w_0573_);
or (w_1465_, w_0699_, w_3511_);
not (w_1385_, w_3255_);
and (w_0943_, w_1879_, w_1329_);
and (w_1014_, w_3510_, w_1767_);
not (w_0000_, in11[6]);
or (w_3098_, w_0906_, w_2647_);
or (w_1796_, w_1787_, w_1105_);
and (w_3006_, in12[0], w_3160_);
and (w_3174_, w_0069_, w_1738_);
or (w_2697_, w_2235_, w_1601_);
or (w_2031_, w_2535_, w_1371_);
or (w_1435_, w_0555_, w_3093_);
and (w_1921_, w_3229_, w_1009_);
not (w_1187_, in2[4]);
or (w_3347_, w_1931_, w_0078_);
or (w_2481_, w_1758_, w_1874_);
and (w_2390_, w_1878_, w_2274_);
and (out15[5], w_1406_, w_0837_);
or (w_2307_, w_0539_, w_2728_);
or (out11[4], w_1610_, w_0757_);
or (w_2061_, w_0705_, w_2256_);
and (w_0747_, w_2204_, w_1528_);
or (w_0082_, w_1317_, w_2097_);
and (w_1041_, in12[1], w_0777_);
and (w_1206_, w_0907_, w_3030_);
and (w_3523_, w_0917_, w_2055_);
or (w_0503_, w_2935_, w_0873_);
or (w_3517_, w_2648_, w_1935_);
and (w_2867_, w_0688_, w_1300_);
and (w_3332_, w_1865_, w_2368_);
not (w_0054_, w_1129_);
or (w_0350_, w_0034_, w_3183_);
and (w_1327_, w_1274_, w_0404_);
or (w_2499_, w_0185_, w_0964_);
and (w_0073_, w_1409_, w_0430_);
or (w_1094_, in9[1], in10[1]);
or (w_2495_, w_0894_, w_1711_);
or (w_2175_, w_2074_, w_1880_);
or (w_3068_, w_2091_, w_0444_);
or (w_1949_, w_0191_, w_2770_);
and (w_1697_, w_0688_, w_2356_);
not (w_1738_, w_2900_);
or (w_3176_, in9[4], in10[4]);
or (out22[7], w_1358_, w_3010_);
and (w_3195_, w_0099_, w_0197_);
not (w_2072_, in9[5]);
or (w_2633_, w_0382_, w_1885_);
and (w_1314_, w_0937_, out13[4]);
not (w_1721_, w_0670_);
and (w_1356_, w_2277_, w_1688_);
or (w_0111_, in11[0], w_1228_);
and (w_3450_, w_3128_, w_0495_);
or (w_0150_, w_2555_, w_2621_);
not (w_1517_, w_1130_);
not (w_2834_, w_2582_);
or (w_2339_, w_2010_, w_1893_);
and (w_2656_, w_3429_, w_0064_);
not (w_0236_, w_1228_);
and (w_3157_, w_0924_, w_1530_);
or (w_1349_, w_1770_, w_3439_);
or (w_1671_, in12[4], w_1678_);
not (w_2855_, w_3276_);
or (w_2859_, w_2345_, w_1800_);
and (w_2590_, w_2049_, w_2132_);
or (w_0706_, in8[0], w_1238_);
and (w_0021_, w_0889_, w_0533_);
and (w_1397_, w_3335_, w_3254_);
and (w_0382_, w_1736_, w_0794_);
and (w_2051_, w_1093_, w_0314_);
and (w_0335_, w_1452_, w_3332_);
and (w_0398_, w_1519_, w_1025_);
not (w_3005_, w_1381_);
and (w_2471_, in11[7], w_1822_);
and (w_3275_, w_1859_, w_1312_);
and (w_2401_, w_1937_, w_1724_);
and (w_0182_, w_2098_, w_2875_);
or (w_2399_, w_0214_, w_2175_);
not (w_1221_, w_2606_);
or (w_0729_, w_2518_, w_2009_);
or (w_2090_, w_2712_, w_1728_);
and (w_3473_, w_2185_, w_1811_);
and (w_1250_, w_1473_, w_2376_);
or (w_2123_, w_2149_, w_0537_);
or (w_3431_, w_2144_, w_2513_);
and (w_0144_, w_1593_, w_1071_);
and (w_1988_, w_3124_, w_0482_);
and (w_3030_, w_1632_, w_1170_);
or (w_0885_, in3[0], w_0328_);
and (w_1982_, w_3074_, w_1394_);
or (w_1298_, in8[1], w_0552_);
not (w_3302_, in13[3]);
not (w_1401_, w_0237_);
and (w_0139_, in8[5], w_1061_);
or (w_0327_, w_2735_, w_2458_);
or (w_1064_, w_2254_, w_1810_);
and (w_2121_, w_1442_, w_0088_);
not (w_0600_, w_2673_);
not (w_2520_, w_3045_);
and (w_0692_, w_3020_, w_0124_);
or (w_1607_, w_2099_, w_1330_);
or (w_2522_, w_3122_, w_0995_);
and (w_0701_, w_2432_, w_2657_);
or (w_1645_, w_1429_, w_0002_);
or (w_0184_, w_1419_, w_1993_);
not (w_0041_, w_2563_);
not (w_0320_, w_0590_);
not (w_0792_, w_2496_);
or (w_0151_, w_3178_, w_2433_);
not (w_2346_, w_2777_);
and (w_0085_, w_1628_, w_2970_);
not (w_3085_, in12[6]);
or (out9[5], w_2268_, w_1681_);
not (w_1555_, in14[0]);
and (w_3255_, w_2014_, w_0201_);
or (w_2293_, w_0113_, w_1999_);
or (w_2700_, w_2924_, w_2662_);
or (w_2507_, w_2639_, w_2342_);
and (w_2223_, in16[0], w_3079_);
or (w_2573_, w_2548_, w_1794_);
and (w_0563_, w_2194_, w_0194_);
or (out16[3], w_1503_, w_2969_);
not (w_2095_, w_2730_);
and (w_3376_, w_0681_, w_0247_);
and (w_1581_, in6[2], in5[1]);
or (w_1494_, w_2598_, w_3124_);
and (w_0211_, w_0322_, w_0016_);
not (w_1945_, w_3443_);
or (out12[0], w_2036_, w_3324_);
and (w_1703_, w_3489_, w_0392_);
and (w_1255_, w_0038_, w_2250_);
or (w_0246_, w_1715_, w_0067_);
and (w_2634_, w_1407_, w_0344_);
or (w_2959_, w_0518_, w_3137_);
not (w_1025_, w_3330_);
and (w_1530_, w_0536_, w_3250_);
and (w_1746_, in1[5], in2[5]);
and (w_3475_, w_0135_, w_2972_);
or (w_0271_, w_0066_, w_2222_);
or (w_0457_, w_2725_, w_0565_);
and (w_0625_, w_1395_, w_3276_);
and (w_2511_, w_1507_, w_0169_);
not (w_2955_, w_3494_);
or (w_1343_, w_0666_, w_1030_);
and (out24[6], w_0560_, w_2155_);
not (w_0493_, w_1936_);
or (w_1271_, w_0099_, w_0197_);
not (w_2243_, in13[2]);
or (w_2962_, w_1056_, w_1537_);
or (w_2423_, w_0456_, w_0501_);
or (w_0377_, w_1628_, w_2970_);
or (out18[3], w_3510_, w_3426_);
or (w_2238_, w_0045_, w_3187_);
and (w_2949_, w_0615_, w_3508_);
or (w_3240_, w_3060_, w_0434_);
and (w_1290_, w_1429_, w_0002_);
or (w_0926_, w_1429_, w_3060_);
and (w_1521_, w_3429_, w_2420_);
or (w_2234_, w_3095_, w_2657_);
and (w_1515_, w_2952_, w_0821_);
and (w_2407_, w_3246_, w_1658_);
or (w_2351_, w_0923_, w_0324_);
not (w_2408_, in14[2]);
not (w_1380_, w_0214_);
and (w_1161_, w_2414_, w_1634_);
and (w_2465_, w_3294_, w_1134_);
not (w_2207_, in3[3]);
and (w_0616_, in9[4], in10[4]);
not (w_1757_, w_3216_);
or (out18[2], w_1393_, w_0217_);
and (w_1684_, w_2991_, w_2004_);
or (w_2086_, w_3516_, w_2678_);
and (w_0577_, w_0990_, w_0773_);
and (w_1708_, w_0963_, w_1424_);
or (w_0008_, w_3203_, w_0018_);
and (w_1883_, w_3330_, w_2669_);
and (w_1463_, w_0991_, w_1428_);
or (w_0286_, w_0471_, w_2052_);
not (w_0448_, w_2803_);
not (w_1539_, w_2511_);
and (w_2777_, w_0900_, w_2748_);
and (w_3087_, w_0482_, w_1336_);
not (w_3296_, w_0157_);
not (w_1855_, w_1464_);
and (w_2996_, w_0906_, w_2647_);
and (w_2967_, w_0161_, w_0504_);
or (w_1809_, in15[6], in16[6]);
or (out21[7], w_0739_, w_0817_);
or (w_2653_, w_0318_, w_0053_);
or (w_2081_, w_1393_, w_0056_);
and (w_2889_, w_1605_, w_2577_);
not (w_3282_, w_1574_);
or (w_2698_, w_1621_, w_0056_);
and (w_3167_, w_2959_, w_2131_);
or (w_0608_, w_1383_, w_0274_);
and (w_3075_, w_1860_, w_3121_);
and (w_2862_, w_1529_, w_0905_);
and (w_2410_, w_2455_, w_1902_);
and (w_1414_, w_0892_, w_0998_);
or (w_1227_, w_1691_, w_2934_);
and (w_2943_, w_1123_, w_1946_);
or (w_1303_, w_2532_, w_1600_);
and (w_2328_, w_2459_, w_2406_);
or (out9[0], w_1772_, w_3418_);
or (out2[5], w_1296_, w_2754_);
or (w_1033_, w_1315_, w_2346_);
or (w_1631_, in13[5], w_3359_);
and (w_2851_, in4[1], w_2327_);
and (w_0670_, in9[5], in10[1]);
and (w_2833_, w_1280_, w_2410_);
not (w_2135_, w_0349_);
and (w_2754_, w_2730_, w_0037_);
and (w_1692_, w_0302_, w_0664_);
or (w_0708_, w_2957_, w_3091_);
or (w_0655_, w_1007_, w_2230_);
not (w_2447_, w_1301_);
not (w_1837_, w_2079_);
and (w_1868_, w_0416_, w_1989_);
and (w_0731_, w_0985_, w_2130_);
or (w_1737_, w_3329_, w_0922_);
or (w_2831_, w_3151_, w_1402_);
or (w_1830_, w_0049_, w_1635_);
or (w_2459_, w_0048_, w_2721_);
not (w_2429_, w_2665_);
and (w_2526_, w_1802_, w_2248_);
or (w_1109_, w_2708_, w_0930_);
or (w_1869_, w_0790_, w_3021_);
and (w_3303_, w_1966_, w_1608_);
or (w_0229_, w_3474_, w_0868_);
or (w_3039_, w_1972_, w_0931_);
and (w_0890_, w_3363_, w_1389_);
or (w_1004_, w_3039_, w_3510_);
or (out18[4], w_0322_, w_2961_);
or (w_0606_, in5[4], w_1659_);
not (w_3124_, w_0804_);
or (w_1674_, w_1981_, w_0713_);
and (w_1600_, w_0921_, w_2404_);
or (w_2432_, w_1697_, w_0949_);
or (w_1415_, w_0769_, w_3382_);
and (w_2852_, w_0450_, w_1344_);
or (w_1381_, w_0034_, w_1174_);
and (w_0592_, w_0379_, w_0628_);
or (w_1427_, in6[5], in5[4]);
or (w_1975_, in15[3], in16[3]);
and (w_2077_, w_3426_, w_2401_);
not (w_2131_, w_1714_);
and (w_1279_, w_2019_, w_2371_);
or (w_2474_, w_0355_, w_0564_);
and (w_3106_, w_2235_, w_1601_);
or (w_2154_, w_2010_, w_0605_);
or (w_0738_, w_0490_, w_3327_);
or (w_1243_, w_1740_, w_0635_);
not (w_2099_, w_3067_);
or (w_1406_, w_3334_, w_1954_);
and (w_0498_, w_0258_, w_3422_);
not (w_1597_, w_0372_);
or (w_1718_, w_1091_, w_3500_);
or (w_0996_, w_2512_, w_1760_);
or (w_1518_, w_1440_, w_2663_);
or (out12[1], w_1795_, w_2030_);
or (w_3407_, w_2918_, w_1054_);
or (w_2577_, w_2893_, w_3127_);
or (w_0855_, w_3492_, w_2526_);
and (w_1457_, w_3452_, w_1912_);
or (w_3043_, w_0076_, w_2188_);
not (w_2694_, w_1521_);
and (w_1257_, w_1110_, w_1492_);
and (w_1228_, w_1292_, w_0364_);
or (w_1820_, w_1097_, w_3326_);
not (w_1442_, w_0550_);
not (w_3022_, w_2094_);
or (w_0886_, w_0707_, w_0597_);
and (w_2063_, w_0803_, w_3486_);
or (w_3149_, w_1746_, w_0847_);
or (w_1896_, w_2371_, w_1320_);
not (w_2854_, w_1758_);
not (w_2882_, in16[7]);
or (w_3365_, out14[3], w_3332_);
or (out13[5], w_1772_, w_3418_);
or (w_2038_, w_1241_, w_2617_);
or (w_2972_, in4[3], w_1205_);
and (w_2654_, w_1949_, w_2820_);
and (w_2279_, w_0441_, w_2607_);
and (w_3398_, w_0790_, w_1969_);
or (w_0481_, w_0461_, w_1490_);
and (w_1351_, w_2506_, w_3036_);
and (w_0777_, w_1013_, w_3485_);
and (out14[3], w_3056_, w_1614_);
or (w_2623_, w_2291_, w_0157_);
or (w_1918_, w_0095_, w_2928_);
or (w_2050_, w_0802_, w_2517_);
or (w_2738_, in9[5], in10[1]);
not (w_0986_, w_1051_);
and (w_2492_, w_0125_, w_3046_);
and (w_2383_, w_2304_, w_0468_);
and (w_1373_, w_2039_, w_0239_);
or (w_0648_, w_1217_, w_3080_);
not (w_0948_, in2[0]);
and (w_1531_, w_2993_, w_1234_);
or (w_0500_, w_0482_, w_1898_);
and (w_2761_, w_0519_, w_3072_);
or (w_3384_, w_0421_, w_0631_);
or (w_1464_, w_2292_, out16[5]);
and (w_1893_, w_3057_, w_2152_);
and (w_2947_, w_0023_, w_2081_);
or (w_0953_, w_0946_, w_0535_);
and (w_1849_, w_2359_, w_2405_);
or (w_0332_, w_0187_, w_0251_);
and (w_3343_, w_3355_, w_2857_);
and (w_0077_, w_0205_, w_1040_);
and (w_0055_, w_0942_, w_0848_);
and (w_3271_, w_0712_, w_2282_);
or (w_1115_, w_2854_, w_0825_);
or (w_2295_, w_0770_, w_1204_);
and (w_3249_, w_2831_, w_0334_);
not (w_2294_, w_1103_);
or (out3[4], w_0958_, w_0891_);
and (out13[1], w_3067_, w_2930_);
or (w_3428_, w_1036_, w_0969_);
and (w_0061_, w_0372_, w_2270_);
and (w_2764_, w_1083_, w_2644_);
or (w_1693_, in16[2], w_1619_);
and (w_2053_, w_3234_, w_2258_);
and (w_1080_, w_1511_, w_2231_);
and (w_0296_, w_2701_, w_1013_);
and (w_2948_, w_1329_, w_0121_);
and (w_1760_, w_1427_, w_1486_);
or (w_2168_, in3[2], w_3303_);
not (w_1797_, w_0208_);
not (w_1801_, w_1818_);
not (w_2120_, w_2790_);
or (w_3394_, w_0877_, w_0525_);
not (w_2206_, w_1166_);
and (w_3349_, w_1714_, w_1383_);
or (w_2735_, w_0798_, w_3106_);
not (w_1665_, w_3308_);
or (w_1749_, w_3012_, w_1957_);
and (w_0714_, w_0214_, w_2175_);
or (w_2017_, w_2451_, w_0899_);
and (w_1346_, in5[4], w_1659_);
or (w_1285_, w_0028_, w_1727_);
or (w_1190_, w_2923_, w_1258_);
not (w_2203_, w_1576_);
or (out20[6], w_1868_, w_0127_);
or (w_0203_, w_1527_, w_1481_);
and (w_2800_, w_1720_, w_1925_);
or (w_1321_, w_1442_, w_0088_);
not (w_2009_, w_2371_);
and (w_0578_, w_2819_, w_1052_);
or (w_0632_, w_2093_, w_3032_);
and (w_1215_, w_3073_, w_3306_);
and (w_3253_, w_0946_, w_0535_);
and (w_3153_, w_2013_, w_3185_);
not (w_0089_, in11[1]);
not (w_2688_, w_0334_);
and (w_1092_, w_0138_, w_0634_);
or (out23[5], w_2085_, w_1821_);
or (w_0494_, w_0045_, w_3361_);
not (w_3337_, w_0109_);
or (w_1491_, w_0000_, w_3256_);
and (w_2752_, w_0094_, w_0327_);
not (w_2510_, w_3105_);
or (w_3212_, w_2814_, w_2122_);
and (w_2370_, w_1522_, w_0289_);
or (w_2318_, in7[2], w_2752_);
or (w_1062_, w_0941_, w_3371_);
or (out10[5], w_1917_, w_3123_);
and (w_0440_, w_0998_, w_1178_);
and (w_3300_, w_0442_, w_2192_);
and (w_2795_, in4[0], w_2994_);
and (w_2079_, in14[7], in13[7]);
or (w_0293_, w_1108_, w_1376_);
and (w_1140_, w_0667_, w_0754_);
or (w_1986_, w_0041_, w_1384_);
and (w_2574_, w_0454_, w_1657_);
and (out22[6], w_0029_, w_2911_);
or (w_2129_, w_1366_, w_2260_);
not (w_2261_, w_2976_);
and (w_1122_, in9[0], in10[0]);
and (w_3155_, w_3213_, w_1073_);
not (w_2548_, w_3108_);
or (w_1934_, w_1155_, w_2855_);
or (w_0553_, w_2796_, w_2159_);
not (w_2472_, w_2649_);
or (w_3361_, w_2572_, w_0763_);
and (w_1831_, w_0904_, w_2606_);
or (w_0044_, w_0487_, w_0158_);
or (w_0038_, w_1110_, w_1492_);
or (w_2676_, w_0889_, w_0533_);
or (w_1101_, w_1679_, out16[1]);
not (w_0118_, in2[2]);
or (w_2946_, w_3168_, w_0967_);
or (out7[5], w_3226_, w_2835_);
or (w_0628_, w_1842_, w_0879_);
and (w_2611_, w_2477_, w_3450_);
or (w_0754_, w_3510_, w_3297_);
not (w_0345_, w_0405_);
and (w_3457_, w_1699_, w_0455_);
or (w_2648_, w_0539_, w_2247_);
or (w_1812_, w_3322_, w_1257_);
or (w_0388_, w_2282_, w_0601_);
and (w_1437_, in4[4], w_0765_);
and (w_0627_, w_1869_, w_1378_);
not (w_3286_, w_3231_);
or (w_0549_, in13[1], w_2127_);
and (w_2479_, in6[5], w_1664_);
or (w_1045_, w_1890_, w_3223_);
and (w_2718_, w_0010_, w_3392_);
and (w_0819_, w_2703_, w_2154_);
and (w_3238_, w_1597_, w_1942_);
and (w_2176_, w_1182_, w_1894_);
and (w_3189_, in4[2], w_1930_);
or (w_3001_, in9[6], in10[2]);
or (w_0474_, in3[3], w_0266_);
or (w_1018_, w_2254_, w_0401_);
and (w_0989_, in14[1], w_2842_);
and (w_2587_, w_0501_, w_2387_);
and (w_1484_, w_2322_, w_0425_);
not (w_2044_, w_1578_);
not (w_0087_, w_3159_);
and (w_2378_, w_0221_, w_3004_);
and (w_0574_, w_0269_, w_3402_);
and (w_1151_, w_1842_, w_3259_);
or (w_2582_, w_1295_, w_0176_);
and (w_1042_, w_1360_, w_0632_);
not (w_3334_, w_2292_);
and (w_3224_, w_1131_, w_1159_);
and (w_2864_, in11[4], w_1287_);
or (w_2705_, w_0461_, w_1752_);
and (w_2604_, w_0441_, w_0361_);
not (w_2384_, w_1996_);
or (w_2606_, in14[7], w_2482_);
or (w_1212_, w_2841_, w_2498_);
and (w_3133_, w_0698_, w_3307_);
and (w_2010_, in1[4], in2[4]);
and (w_2052_, w_2415_, w_2478_);
and (w_1177_, w_1466_, w_0214_);
and (w_1012_, w_0661_, w_1310_);
or (w_3522_, in11[6], w_1237_);
and (w_0412_, w_2701_, w_3230_);
and (w_1231_, w_0601_, w_0710_);
and (w_1069_, in9[5], in10[5]);
and (w_2564_, w_2648_, w_1935_);
not (w_1804_, w_2231_);
and (w_0717_, w_2813_, w_0792_);
and (w_0573_, w_3188_, w_2375_);
and (w_0674_, w_2614_, w_1324_);
or (w_1498_, w_0417_, w_2949_);
and (w_1507_, w_0940_, w_3340_);
and (w_2668_, w_3275_, w_1796_);
or (w_0726_, w_0851_, w_2966_);
and (w_2434_, w_0735_, w_1444_);
or (w_1044_, w_3248_, w_2913_);
and (w_1980_, w_2639_, w_2342_);
or (w_0270_, w_3225_, w_1775_);
and (w_3205_, in12[6], w_3061_);
and (w_1947_, w_1823_, w_1254_);
and (w_2242_, w_1258_, w_2961_);
and (w_2650_, in6[4], w_0526_);
or (w_3503_, w_0601_, w_3081_);
or (w_0396_, w_1961_, w_2782_);
or (w_2868_, w_0144_, w_2311_);
and (w_1220_, w_3101_, w_1032_);
or (w_1723_, w_2618_, w_2019_);
or (w_2911_, w_2463_, w_0592_);
or (w_1142_, in6[2], w_0440_);
and (w_0643_, w_0655_, w_1168_);
not (w_2286_, w_0507_);
or (w_1458_, in15[6], w_2361_);
and (w_0053_, w_2345_, w_1800_);
or (w_2155_, out14[6], w_2672_);
and (w_2193_, in3[0], w_2940_);
and (w_2513_, w_0008_, w_0606_);
not (w_2450_, w_0044_);
or (w_2682_, w_2452_, w_0278_);
or (w_0084_, w_0804_, w_1150_);
and (w_0694_, in15[6], w_2361_);
or (w_0297_, w_3454_, w_0588_);
or (w_0589_, w_3503_, w_0222_);
and (w_0489_, w_2974_, w_1176_);
and (w_1968_, w_3454_, w_0588_);
or (w_2641_, w_2402_, w_1704_);
and (w_3014_, w_1986_, w_1438_);
not (w_1201_, w_0043_);
or (w_1626_, w_0689_, out16[0]);
or (w_1989_, w_3369_, w_1078_);
and (w_3320_, w_1477_, w_0513_);
or (w_3242_, w_3316_, w_2608_);
or (w_0279_, w_1144_, w_0318_);
not (w_1422_, w_2727_);
not (w_0688_, w_2618_);
or (w_0083_, w_3406_, w_2161_);
and (w_2483_, w_0443_, w_0976_);
and (out7[1], w_1152_, w_2891_);
or (w_1431_, w_0417_, w_0462_);
or (w_0920_, out14[2], w_1949_);
and (w_2780_, w_2409_, w_3506_);
and (w_2965_, w_2146_, w_0306_);
or (w_0187_, w_0751_, w_1471_);
not (w_2114_, w_3026_);
or (w_1676_, w_2199_, w_1546_);
and (w_2274_, w_1522_, w_2486_);
not (w_1441_, w_2687_);
and (out9[1], w_2649_, w_1701_);
or (w_2353_, w_1529_, w_0905_);
or (out12[5], w_0308_, w_0701_);
or (w_2584_, w_1415_, w_0478_);
and (w_1087_, w_0942_, w_1549_);
or (w_1132_, in1[4], in2[4]);
and (w_1818_, w_1552_, w_1158_);
or (w_1902_, in8[3], w_2145_);
and (w_0417_, in15[4], in16[4]);
not (w_2670_, w_1526_);
or (w_2054_, w_0438_, w_1163_);
and (w_3257_, w_2111_, w_2885_);
or (w_1932_, w_0866_, w_1241_);
or (w_2936_, w_0840_, w_2424_);
or (w_0304_, in14[5], w_2777_);
and (w_1747_, w_1864_, w_2021_);
or (w_2897_, w_3192_, w_1306_);
or (w_1233_, w_1119_, w_0516_);
or (w_1260_, w_2034_, w_0595_);
or (w_0225_, w_2072_, w_2302_);
and (w_2397_, w_1089_, w_0816_);
or (w_0497_, w_2437_, w_3425_);
or (w_0306_, w_2411_, w_3449_);
or (w_1808_, w_3398_, w_0402_);
and (out6[4], w_1842_, w_2803_);
or (w_0900_, w_1824_, w_2262_);
and (w_0070_, w_0657_, w_2791_);
or (w_1907_, w_1789_, w_1387_);
or (w_2320_, w_0815_, w_2844_);
or (w_0072_, in12[0], w_2745_);
or (w_1513_, w_3105_, w_1022_);
or (w_2536_, w_3456_, w_0052_);
not (w_0245_, w_3479_);
and (w_1107_, w_0653_, w_1403_);
or (w_3086_, w_2808_, w_3338_);
or (w_2259_, w_0449_, w_3300_);
or (w_2305_, w_2321_, w_1862_);
and (w_1481_, w_1717_, w_3119_);
and (w_1770_, w_0646_, w_2816_);
or (w_3110_, w_0209_, w_0369_);
and (w_0458_, w_1200_, w_2673_);
not (w_1426_, w_2491_);
or (w_2980_, w_1053_, w_1934_);
or (w_3499_, w_2921_, w_0984_);
not (w_1623_, w_1408_);
and (w_2411_, in6[2], w_0440_);
and (w_0713_, w_2761_, w_2597_);
and (w_2358_, w_0790_, w_3385_);
or (w_1724_, w_3165_, w_0353_);
and (w_0564_, w_0671_, w_2518_);
and (w_2957_, w_3034_, w_1566_);
not (w_1420_, in4[0]);
not (w_1987_, w_0408_);
not (w_1000_, w_1345_);
or (w_2149_, w_2881_, w_1332_);
or (w_3269_, w_0216_, w_2880_);
or (w_3115_, in14[4], w_3466_);
not (w_3482_, w_0028_);
and (w_0828_, w_0733_, w_2679_);
or (w_1864_, w_2295_, w_3512_);
and (w_2810_, w_2007_, w_1591_);
not (w_2926_, w_0125_);
and (w_3026_, w_3434_, w_0801_);
and (w_1209_, in12[5], w_0740_);
and (w_0287_, out14[6], w_2672_);
or (w_2610_, in7[3], w_3257_);
and (w_0758_, w_0317_, w_3113_);
not (w_2721_, w_3158_);
or (w_1519_, w_2066_, w_3271_);
or (w_3237_, w_1871_, w_1018_);
or (w_0202_, in6[3], in5[2]);
and (w_0027_, w_0689_, out16[0]);
and (w_1691_, in8[4], w_2751_);
or (w_3280_, w_1662_, w_0590_);
not (w_3011_, w_3144_);
not (w_0551_, w_0609_);
not (w_1582_, w_0947_);
and (w_3313_, w_0790_, w_2019_);
and (w_3031_, w_3405_, w_2303_);
or (out23[7], w_2164_, w_2082_);
and (w_3160_, w_1147_, w_2746_);
and (w_2770_, w_3328_, w_2388_);
and (w_0291_, w_0263_, w_3241_);
and (w_0576_, w_0889_, w_2076_);
not (w_2141_, w_3175_);
or (w_1405_, w_2185_, w_1811_);
or (w_0997_, w_2202_, w_0368_);
or (w_1146_, w_0138_, w_0634_);
or (w_3357_, w_2847_, w_1267_);
or (w_2270_, w_2839_, w_2384_);
and (w_2835_, w_1963_, w_0627_);
or (w_0312_, w_1380_, w_1242_);
or (out11[2], w_2538_, w_0674_);
not (w_2182_, w_1458_);
not (w_2525_, w_0304_);
or (w_0641_, w_2194_, w_2438_);
or (w_1291_, w_1877_, w_1761_);
or (w_1068_, w_0294_, w_1106_);
not (w_3051_, w_0873_);
and (w_2458_, w_0272_, w_1142_);
and (w_0784_, w_2819_, w_2332_);
and (w_2994_, w_1740_, w_0384_);
or (out10[3], w_0861_, w_0027_);
or (out19[6], w_1246_, w_0248_);
and (w_1992_, w_3325_, w_3020_);
and (w_2247_, w_2340_, w_3521_);
and (w_0075_, w_2115_, w_2058_);
and (w_0356_, w_1173_, w_1779_);
not (w_0956_, in9[0]);
and (w_3227_, w_0120_, w_0103_);
and (w_1270_, w_1463_, out16[6]);
and (w_0585_, w_1198_, w_0645_);
not (w_0536_, w_2611_);
or (w_2872_, w_3379_, w_1840_);
or (w_0399_, w_0296_, w_1392_);
and (w_1493_, w_0923_, w_0324_);
and (w_0265_, w_1756_, w_3082_);
and (w_2043_, w_0774_, w_1594_);
or (w_0379_, w_0221_, w_2428_);
or (w_0058_, w_0488_, w_3249_);
not (w_2715_, w_0492_);
or (w_2023_, w_2724_, w_3208_);
not (w_2227_, w_2501_);
not (w_1798_, w_3132_);
or (out23[0], w_1140_, w_1289_);
and (w_3464_, w_3325_, w_2734_);
or (w_2255_, w_2515_, w_1667_);
or (w_3485_, w_0128_, w_0412_);
and (w_2837_, w_2064_, w_2504_);
and (w_1634_, w_1278_, w_0542_);
and (w_0156_, out13[6], w_3418_);
and (w_2301_, w_1827_, w_1082_);
and (w_3342_, w_0501_, w_0173_);
not (w_3409_, w_0303_);
or (w_2442_, w_0774_, w_1594_);
or (w_2025_, w_2365_, w_3462_);
and (w_0770_, w_2017_, w_0791_);
or (w_1253_, w_3034_, w_3528_);
or (w_1364_, w_0870_, w_2688_);
or (w_0140_, w_3492_, w_1329_);
and (w_0496_, w_3510_, out13[0]);
not (w_1566_, w_1531_);
and (w_1425_, w_1081_, w_0980_);
and (w_0710_, w_2849_, w_3393_);
or (w_0937_, w_0534_, w_0761_);
or (w_2981_, w_0671_, w_0217_);
and (w_3141_, w_3218_, w_0781_);
not (w_2348_, w_1547_);
or (w_2150_, w_0989_, w_2015_);
and (w_2559_, in14[5], w_2107_);
or (w_0779_, in1[5], in2[5]);
or (w_1939_, w_0671_, w_2518_);
not (w_3088_, w_2600_);
not (w_2211_, w_2122_);
and (w_3392_, w_0749_, w_2032_);
and (w_0217_, w_0547_, w_2583_);
not (w_0994_, w_0826_);
and (w_1735_, w_3242_, w_2836_);
or (w_0637_, w_1926_, w_2862_);
not (w_3256_, w_1237_);
or (w_3162_, w_2938_, w_1974_);
or (w_3246_, w_0506_, w_0315_);
and (w_1941_, w_0851_, w_2966_);
not (w_0734_, w_1308_);
or (w_3393_, w_1535_, w_0271_);
and (w_1688_, w_2661_, w_1578_);
or (w_1395_, w_3041_, w_0593_);
or (w_1275_, w_2244_, w_3051_);
or (w_2791_, w_2922_, w_2391_);
and (w_0883_, w_0617_, w_3459_);
and (w_0804_, w_0031_, w_2045_);
not (w_2382_, w_1031_);
and (w_0278_, w_3316_, w_0330_);
or (w_2409_, w_1024_, w_1580_);
and (w_1618_, w_1068_, w_0012_);
or (w_1615_, w_1102_, w_1143_);
not (w_0437_, w_2404_);
or (w_3117_, w_1393_, w_0671_);
and (w_2089_, w_1996_, w_0405_);
not (w_2310_, w_0209_);
and (w_3024_, w_0802_, w_3263_);
not (w_0669_, w_1095_);
or (out16[4], w_1223_, w_2242_);
or (w_2543_, w_3247_, w_2654_);
not (w_2873_, in3[0]);
and (w_3471_, w_1707_, w_3432_);
or (w_0980_, w_1810_, w_1154_);
or (w_2239_, w_3275_, w_1796_);
or (w_1856_, w_1209_, w_0672_);
or (w_0366_, w_3328_, w_2388_);
and (w_0526_, w_2507_, w_3431_);
and (w_2707_, w_1211_, w_2633_);
and (w_1400_, w_1174_, w_2586_);
not (w_0502_, w_3056_);
or (w_1017_, w_2175_, w_1030_);
not (w_0904_, w_2982_);
or (w_1861_, in14[7], in13[7]);
or (w_0266_, w_2689_, w_2542_);
or (w_2169_, w_3037_, w_0298_);
and (w_2022_, w_2292_, out16[5]);
and (w_2316_, w_2505_, w_1631_);
not (w_2826_, w_1001_);
and (w_2696_, w_1598_, w_1484_);
or (w_0863_, w_3034_, w_1566_);
and (w_1836_, in14[4], in13[4]);
or (w_2692_, w_0322_, w_0237_);
and (w_2556_, w_1071_, w_0721_);
or (w_1440_, w_3505_, w_2893_);
or (w_0867_, w_1616_, w_3330_);
or (w_3077_, w_0599_, w_0489_);
not (w_0051_, w_2488_);
or (w_2684_, w_3492_, w_0512_);
and (w_3016_, w_0774_, w_1809_);
or (w_2069_, w_1971_, w_0299_);
not (w_3436_, w_2839_);
and (w_1117_, w_3497_, w_0073_);
or (w_2585_, w_2467_, w_0955_);
and (w_1061_, w_0996_, w_2977_);
and (w_2365_, w_3424_, w_3416_);
not (w_1957_, w_3346_);
not (w_0164_, w_2678_);
or (w_0888_, w_1401_, w_0844_);
or (w_0046_, w_2839_, w_2089_);
or (w_2603_, w_1273_, w_0473_);
not (w_0846_, w_2392_);
not (w_1111_, in16[4]);
and (w_1974_, w_3172_, w_3386_);
or (w_0326_, w_2046_, w_3215_);
or (w_2026_, w_1883_, w_1282_);
and (w_3070_, in8[3], w_2145_);
not (w_2763_, w_3023_);
not (w_3495_, w_1678_);
or (w_3147_, w_3426_, w_2401_);
and (w_0219_, w_0802_, w_0064_);
or (w_0430_, w_0322_, w_0016_);
or (w_3177_, w_2881_, w_1039_);
and (w_2116_, w_1240_, w_2824_);
and (w_1772_, w_0790_, w_3352_);
and (w_0301_, in12[2], w_0409_);
or (w_3295_, w_0007_, w_0210_);
or (w_2322_, w_2243_, w_1577_);
not (w_2414_, in11[7]);
or (w_0562_, w_2068_, w_2614_);
or (w_0968_, w_1118_, w_0766_);
and (w_3204_, w_2959_, w_0281_);
not (w_1074_, w_1643_);
not (w_1119_, w_1463_);
and (w_0009_, w_3472_, w_1937_);
and (w_0868_, w_1857_, w_1185_);
or (w_2973_, w_1612_, w_0160_);
or (w_1424_, w_1828_, w_0978_);
and (w_0092_, w_2508_, w_0926_);
and (w_3251_, w_2840_, w_3296_);
and (out16[7], w_2035_, w_1469_);
or (w_3472_, w_1452_, w_3332_);
and (w_1951_, w_2261_, w_2020_);
or (w_1085_, w_2792_, w_3476_);
or (w_0619_, w_0804_, w_0421_);
or (w_2885_, w_0653_, w_1403_);
and (w_3494_, w_2062_, w_2495_);
or (out19[1], w_2959_, w_1637_);
and (w_2030_, w_2270_, w_1734_);
or (w_1908_, w_0331_, w_2037_);
and (w_1348_, w_2690_, w_0803_);
or (w_1392_, w_3390_, w_0359_);
and (w_2939_, w_0963_, w_1977_);
and (w_1594_, w_1556_, w_1809_);
or (w_1367_, in4[3], w_1042_);
or (w_1362_, w_1623_, w_2392_);
or (w_0677_, w_1648_, w_1249_);
and (w_1365_, w_2518_, w_1737_);
and (w_2804_, w_3264_, w_2301_);
and (w_3216_, out10[0], w_2485_);
and (w_0927_, in8[2], w_1851_);
and (w_0541_, w_2415_, w_1842_);
not (w_2074_, w_0928_);
not (w_1870_, in9[4]);
and (w_3371_, w_1275_, w_3277_);
or (w_0330_, w_0476_, w_0226_);
or (w_1251_, w_0910_, w_2900_);
and (w_3308_, in12[7], w_2651_);
or (w_1232_, w_0826_, w_3167_);
not (w_3341_, w_1727_);
not (w_1528_, w_2768_);
or (w_0023_, w_0802_, w_3263_);
or (w_0034_, w_0782_, w_1919_);
not (w_0482_, w_3426_);
not (w_1736_, w_2712_);
and (w_2745_, w_0982_, w_0111_);
and (w_2376_, w_0742_, w_0280_);
and (w_1159_, w_1958_, w_0391_);
not (w_2268_, w_1956_);
and (w_1821_, w_0209_, w_0764_);
and (w_2828_, w_2442_, w_3455_);
and (w_1983_, w_2828_, w_1138_);
or (w_0110_, w_3170_, w_1596_);
not (w_1673_, w_0790_);
and (out22[4], w_3086_, w_3499_);
and (w_0499_, in15[0], w_0509_);
not (w_1305_, w_0954_);
and (w_0579_, w_0496_, w_0014_);
or (w_2952_, w_2922_, w_2830_);
and (out13[0], w_0354_, w_2354_);
or (w_3245_, w_3155_, w_1990_);
or (w_0284_, w_2210_, w_1505_);
or (w_0113_, w_2614_, w_0485_);
or (w_1658_, in12[2], w_1461_);
and (w_2457_, in7[4], w_2229_);
and (w_3328_, w_0232_, w_2715_);
and (w_2922_, w_3039_, w_3510_);
and (w_0128_, in11[0], w_1228_);
and (w_1043_, w_0074_, w_0130_);
and (w_0672_, w_0814_, w_2430_);
and (w_3175_, w_0789_, w_2737_);
or (w_0289_, w_0546_, w_1889_);
or (w_3219_, in8[4], w_3184_);
and (w_0238_, w_3248_, w_2913_);
not (w_2579_, in5[3]);
and (w_2183_, w_0839_, w_2432_);
or (w_3486_, w_1398_, w_0575_);
or (w_2117_, w_1301_, w_0256_);
and (w_0318_, w_2285_, w_3099_);
not (w_1791_, w_3269_);
and (w_0461_, in16[2], w_1619_);
not (w_0381_, w_0740_);
and (w_0793_, w_2974_, w_0581_);
or (w_3416_, w_1067_, w_0172_);
and (w_0476_, in11[5], w_1984_);
and (w_1654_, w_2843_, w_0859_);
or (w_1429_, w_2166_, w_1510_);
or (w_1640_, w_2963_, w_1164_);
not (w_1281_, w_0468_);
and (w_1944_, w_2445_, w_0481_);
not (w_1621_, w_2580_);
and (w_3274_, w_2985_, w_2712_);
and (w_1744_, w_2795_, w_3464_);
and (w_1940_, w_3211_, w_1362_);
or (w_1158_, w_0654_, w_2271_);
or (w_0837_, w_2292_, w_0968_);
or (w_2644_, w_0522_, w_1831_);
and (w_2119_, w_0501_, w_0482_);
and (w_1675_, w_2742_, w_0829_);
and (w_0443_, w_0500_, w_3147_);
or (w_2349_, w_1509_, w_2549_);
and (out14[2], w_1907_, w_3354_);
or (w_0973_, in14[0], in13[0]);
or (w_0386_, w_3482_, w_3341_);
not (w_3037_, w_3186_);
or (w_1826_, w_0788_, w_0254_);
and (w_1118_, w_1320_, w_1714_);
or (w_2180_, w_1968_, w_2702_);
not (w_1325_, w_2362_);
or (w_2424_, w_0524_, w_0131_);
and (w_0401_, w_0617_, w_1055_);
and (w_0197_, w_2727_, w_0704_);
and (w_2986_, w_2499_, w_1733_);
and (w_0955_, w_0553_, w_2041_);
and (w_1468_, w_0388_, w_2551_);
not (w_0561_, w_1513_);
or (w_2404_, in12[2], w_0409_);
not (w_1199_, w_1677_);
not (w_1508_, w_2597_);
or (w_0395_, w_2591_, w_0997_);
or (w_1476_, w_1552_, w_2271_);
and (w_0178_, in11[3], w_0643_);
or (w_2887_, in14[1], w_2842_);
or (w_1411_, w_3021_, w_1124_);
not (w_3042_, w_0093_);
or (w_2398_, w_2640_, w_2587_);
or (w_2652_, w_1026_, w_0557_);
or (w_2506_, w_3494_, w_2959_);
and (out7[0], w_0947_, w_2280_);
or (w_0375_, w_0644_, w_0959_);
not (w_0993_, w_1278_);
not (w_1226_, w_3523_);
or (w_2786_, w_0415_, w_0703_);
and (w_0965_, w_2241_, w_3298_);
or (w_2561_, w_2209_, w_3523_);
and (w_3388_, w_2153_, w_3105_);
and (w_1136_, w_3203_, w_0018_);
or (w_1379_, w_0781_, w_3426_);
and (w_0324_, w_0778_, w_1299_);
not (w_3062_, w_2309_);
and (w_3082_, w_2550_, w_2308_);
and (w_1252_, w_2207_, w_0333_);
and (w_1247_, w_0527_, w_3251_);
not (w_0903_, w_3511_);
or (out8[5], w_0785_, w_2389_);
and (w_2392_, w_2371_, w_1022_);
or (w_2343_, w_2223_, w_3009_);
and (w_2356_, w_1265_, w_3076_);
and (w_2373_, w_2729_, w_2453_);
or (w_2992_, w_0284_, w_0100_);
and (w_0343_, in8[1], w_3233_);
not (w_1081_, in8[2]);
or (w_0198_, w_1788_, w_2762_);
and (w_0761_, w_0252_, w_2805_);
not (w_1642_, in10[4]);
and (w_3414_, w_0618_, w_2502_);
not (w_0485_, w_0760_);
not (w_0506_, in12[2]);
or (w_1152_, w_0947_, w_2075_);
and (w_2744_, w_2973_, w_0231_);
or (w_1546_, w_0683_, w_2546_);
or (w_1169_, w_3066_, w_3054_);
not (w_0339_, in1[0]);
not (w_2068_, w_0271_);
and (w_1482_, w_1395_, w_2980_);
and (w_2174_, w_1150_, w_0671_);
and (w_0409_, w_0399_, w_2123_);
not (w_0699_, w_3001_);
and (w_2659_, w_1651_, w_3421_);
and (w_2599_, w_1719_, w_1535_);
or (w_1423_, w_0421_, w_1895_);
and (w_2782_, w_3186_, w_2011_);
or (w_0311_, in14[3], in13[3]);
or (w_1030_, w_0115_, w_3447_);
or (w_2870_, w_0865_, w_1245_);
and (w_0142_, w_2128_, w_2956_);
or (w_0160_, w_0346_, w_3000_);
not (w_2466_, w_1160_);
and (w_0338_, w_1320_, w_0659_);
or (w_1408_, w_2371_, w_1022_);
and (w_2219_, w_1408_, w_0846_);
or (w_1553_, w_2408_, w_1572_);
not (w_0022_, w_0754_);
and (w_2240_, w_0421_, w_2009_);
and (w_1471_, w_2618_, w_2518_);
or (w_3380_, w_3211_, w_1362_);
or (w_3277_, w_3236_, w_0873_);
not (w_1875_, w_1927_);
and (w_0331_, w_2566_, w_0859_);
or (w_0255_, w_0340_, w_0165_);
and (w_2956_, w_0063_, w_1782_);
and (w_2394_, w_2025_, w_2351_);
or (w_0020_, w_3377_, w_1825_);
and (w_3340_, w_0394_, w_2876_);
and (w_0546_, w_2129_, w_2111_);
not (w_0571_, w_1371_);
not (w_0548_, w_2177_);
or (w_2204_, w_1463_, w_2767_);
and (w_2202_, in13[7], w_3038_);
or (w_0657_, w_0253_, w_3322_);
or (out20[5], w_2469_, w_2547_);
and (w_1979_, w_0970_, w_2112_);
or (w_2944_, w_1866_, w_0246_);
not (w_1098_, w_0957_);
or (w_3470_, w_0039_, w_3265_);
and (w_0467_, w_1666_, w_3050_);
not (w_0748_, w_0857_);
or (w_3476_, w_1595_, w_3214_);
and (w_2827_, w_2419_, w_0114_);
or (w_0241_, w_0252_, out13[3]);
or (w_1690_, in3[5], w_1531_);
or (w_0610_, w_2069_, w_0517_);
or (w_2273_, w_2722_, w_1872_);
or (w_2363_, w_0387_, w_2686_);
not (w_0102_, w_2593_);
or (w_1653_, w_2627_, w_2632_);
and (w_0582_, in16[5], w_0090_);
or (w_2811_, w_1991_, w_2255_);
or (w_2635_, w_2358_, w_2719_);
and (w_1596_, w_2131_, w_2672_);
and (w_2171_, w_0612_, w_2374_);
and (w_1871_, w_2363_, w_2054_);
or (w_0392_, w_1707_, w_3432_);
or (w_0522_, w_1155_, w_0307_);
and (w_1571_, w_2297_, w_3448_);
and (w_1195_, w_2101_, w_0890_);
and (w_3453_, w_0214_, w_2803_);
not (w_0453_, w_1961_);
or (w_0629_, w_1386_, w_0348_);
and (w_2988_, w_0449_, w_3300_);
and (w_1217_, w_0836_, w_0863_);
and (out1[0], w_0354_, w_2354_);
or (w_1312_, in5[3], w_3460_);
or (w_2248_, w_0937_, out13[4]);
and (w_2091_, w_0671_, w_0217_);
and (w_3125_, w_1262_, w_1820_);
or (w_1651_, w_3429_, w_0064_);
and (w_0776_, w_0608_, w_3240_);
and (w_2208_, w_2017_, w_1646_);
or (w_0712_, w_3401_, w_0040_);
or (w_1506_, w_1308_, w_2317_);
or (w_1575_, w_2305_, w_2298_);
or (w_2619_, w_0446_, w_0579_);
and (w_0307_, w_3295_, w_0625_);
or (w_2539_, w_2471_, w_1019_);
and (w_2544_, in4[5], w_2945_);
not (w_1901_, w_0572_);
or (w_1806_, w_2266_, w_2314_);
not (w_1514_, w_0092_);
and (w_3107_, w_3001_, w_0903_);
or (w_2249_, w_0985_, w_2130_);
or (w_0639_, w_2726_, w_3028_);
and (w_2709_, w_3445_, w_3094_);
or (w_2533_, w_2034_, w_2065_);
and (w_0067_, in14[0], in13[0]);
and (w_1359_, in1[3], in2[3]);
and (w_0492_, w_1174_, w_0064_);
and (w_0376_, w_3406_, w_2161_);
not (w_0477_, in13[6]);
and (w_0196_, w_0082_, w_0072_);
and (w_3427_, w_2316_, w_0293_);
or (w_0093_, w_0034_, w_2961_);
not (w_1850_, w_0183_);
or (w_1123_, w_3367_, w_2047_);
not (w_2849_, w_1586_);
or (w_1999_, w_1668_, w_1413_);
and (w_2919_, w_2474_, w_1750_);
or (w_2236_, w_0598_, w_2211_);
or (w_0933_, w_2618_, w_2518_);
and (w_1267_, w_1673_, w_1025_);
and (out14[0], w_3503_, w_3017_);
or (w_1120_, w_3013_, w_2557_);
and (w_1054_, w_0970_, w_0902_);
or (w_0814_, w_0410_, w_2950_);
or (w_2433_, w_0871_, w_3409_);
not (w_2289_, w_3155_);
and (w_1417_, w_1849_, out16[7]);
or (w_0358_, w_2386_, w_0611_);
and (w_0852_, w_2895_, w_1174_);
or (w_2875_, w_2421_, w_1005_);
and (w_1833_, w_0228_, w_1121_);
and (w_2877_, w_2870_, w_3434_);
not (w_2425_, w_3513_);
or (w_2509_, w_1091_, w_2638_);
or (w_1657_, in4[1], w_1732_);
and (w_3047_, w_3262_, w_1764_);
and (w_1289_, w_0877_, w_0022_);
not (w_1781_, w_1213_);
and (w_1421_, w_0387_, w_2686_);
or (w_1584_, w_3526_, w_1065_);
or (w_2158_, w_2197_, w_1064_);
not (w_3445_, in8[4]);
not (w_0932_, w_0129_);
not (w_2691_, w_0046_);
and (w_0170_, w_3526_, w_1065_);
not (w_2209_, w_0962_);
and (w_1960_, w_2307_, w_1351_);
and (w_0936_, w_1539_, w_3003_);
not (w_0807_, w_3390_);
or (w_1473_, w_3168_, w_0423_);
or (w_2111_, w_0123_, w_0270_);
and (w_3348_, w_0241_, w_1256_);
and (w_3377_, w_3494_, w_0935_);
or (w_2995_, w_0895_, w_1259_);
or (w_3120_, w_2827_, w_0066_);
and (w_0352_, w_1242_, w_1817_);
or (w_1185_, w_0781_, w_3348_);
or (w_1432_, w_0940_, w_3340_);
or (w_1661_, w_2667_, w_0860_);
or (w_1709_, w_0798_, w_0737_);
not (w_0450_, w_2581_);
or (out20[1], w_1970_, w_1695_);
not (w_3179_, in15[3]);
or (w_1547_, w_1246_, w_3081_);
and (w_1479_, w_1393_, w_1329_);
not (w_2470_, w_1036_);
and (w_1554_, out15[0], w_2225_);
or (w_0581_, w_2895_, w_1174_);
not (w_2360_, w_0491_);
or (w_1756_, w_0796_, w_3401_);
or (w_1728_, w_2590_, w_0177_);
and (out17[5], w_0790_, w_1519_);
or (w_0942_, w_1356_, w_1349_);
or (out12[3], w_2022_, w_1855_);
and (w_0797_, w_3358_, w_0832_);
and (w_0513_, w_2723_, w_1186_);
and (w_0103_, w_0263_, w_2605_);
or (w_3373_, out10[0], w_2485_);
and (w_0317_, w_0698_, w_1966_);
not (w_2789_, w_1451_);
or (w_1477_, w_0870_, w_2975_);
or (w_2102_, w_1195_, w_2541_);
and (w_2999_, w_3036_, w_1316_);
and (w_1559_, w_1479_, w_2190_);
and (w_2106_, w_0264_, w_0186_);
or (w_1297_, w_1150_, w_0671_);
and (w_3207_, w_0322_, w_3248_);
or (w_1916_, w_2348_, w_3171_);
and (w_3265_, w_0804_, w_1150_);
and (out24[5], w_0843_, w_2350_);
not (w_2524_, w_0067_);
and (w_2164_, w_1218_, w_1513_);
or (w_0635_, w_2552_, w_0563_);
or (w_2241_, w_1292_, w_1765_);
and (w_0049_, w_1166_, w_0148_);
not (w_2210_, w_1423_);
or (w_2148_, w_3497_, w_3105_);
or (w_2797_, w_3417_, w_2861_);
and (w_1993_, w_0255_, w_3144_);
and (w_1179_, w_2223_, w_3255_);
not (w_1149_, in11[0]);
or (w_3400_, w_2460_, w_3360_);
and (out21[4], w_0065_, w_0709_);
and (w_2321_, w_3021_, w_1124_);
not (w_1512_, w_3496_);
or (w_1829_, w_2012_, w_0759_);
and (w_1704_, w_2363_, w_1086_);
not (w_2075_, w_1561_);
and (w_3034_, w_2061_, w_1264_);
or (out3[1], w_0835_, w_1819_);
or (w_1698_, w_2366_, w_1781_);
not (w_0715_, w_3072_);
not (w_2142_, w_2170_);
or (w_0580_, w_0104_, w_3495_);
and (w_0491_, w_1607_, out13[2]);
and (w_0030_, w_0291_, w_1685_);
and (w_0552_, w_2054_, w_2641_);
not (w_0516_, w_0234_);
and (w_3395_, w_3293_, w_1020_);
not (w_1799_, in2[3]);
or (w_2381_, w_2336_, w_2079_);
or (w_3462_, w_1670_, w_3458_);
not (w_2096_, in12[5]);
and (w_3184_, w_1271_, w_1502_);
not (w_0001_, w_0187_);
not (w_1378_, w_1143_);
or (w_2032_, in5[1], w_0692_);
and (w_1160_, w_0416_, w_3222_);
and (w_1145_, w_3416_, w_0091_);
and (w_3146_, w_2193_, w_2053_);
or (w_0565_, w_0410_, w_0189_);
and (w_3465_, in13[2], w_1807_);
or (out16[2], w_0636_, w_1500_);
or (w_1852_, w_3057_, w_2152_);
and (w_2822_, w_1636_, w_2278_);
not (w_0525_, w_1343_);
and (w_0603_, w_1028_, w_0780_);
or (w_0787_, w_2335_, w_1255_);
and (w_1342_, w_0804_, w_0421_);
and (w_0439_, w_2870_, w_3115_);
and (out4[1], w_0321_, w_1916_);
and (w_3064_, w_1198_, w_3383_);
and (w_0935_, w_0311_, w_0532_);
or (w_3419_, w_3231_, w_0129_);
and (w_1814_, w_1875_, w_2786_);
or (w_3035_, w_0181_, w_1457_);
not (w_1792_, w_2535_);
and (w_0826_, w_0322_, w_1714_);
and (w_3079_, w_2613_, w_1928_);
or (w_0972_, w_2457_, w_1063_);
or (out19[7], w_0187_, w_2510_);
and (w_0410_, in12[4], w_1678_);
and (w_3263_, w_2104_, w_3437_);
and (w_1237_, w_3062_, w_0977_);
and (w_2391_, w_2282_, w_0601_);
and (w_2190_, w_1242_, w_3248_);
not (w_0341_, w_3153_);
and (w_2201_, w_3074_, w_2887_);
or (w_2625_, in15[4], in16[4]);
not (w_1603_, w_2744_);
not (w_3201_, w_0302_);
not (w_0862_, w_2883_);
not (w_1497_, w_3307_);
not (w_2186_, w_2246_);
and (w_1817_, w_0626_, w_1297_);
and (w_1616_, w_0084_, w_2189_);
not (w_1954_, w_0968_);
not (w_0117_, w_0461_);
or (w_0120_, w_2938_, w_1206_);
not (w_0601_, w_3510_);
and (w_1562_, w_2535_, w_1371_);
or (w_2757_, w_0945_, w_2216_);
or (w_1551_, w_2877_, w_2540_);
or (w_0569_, w_0669_, w_1535_);
and (w_2726_, w_0804_, w_3426_);
or (w_2857_, w_3283_, w_2946_);
and (w_1105_, w_0531_, w_2252_);
and (w_1048_, w_2263_, w_2909_);
or (out13[6], w_0913_, w_0235_);
or (w_2562_, w_0887_, w_0594_);
and (w_2034_, w_1737_, w_0237_);
and (w_1552_, w_1175_, w_2983_);
and (w_2065_, w_2853_, w_2352_);
and (w_3054_, w_0506_, w_0315_);
not (w_0099_, in7[3]);
and (w_0794_, w_1729_, w_0101_);
or (w_0201_, in16[1], w_0208_);
and (w_0333_, w_0378_, w_3520_);
and (w_0915_, w_0697_, w_2024_);
or (w_2143_, w_1598_, w_1484_);
and (w_1337_, w_2831_, w_0207_);
or (w_1079_, w_1235_, w_1627_);
or (w_0774_, w_1097_, w_0192_);
and (w_0799_, w_2234_, w_1112_);
or (out3[0], w_0316_, w_0465_);
and (w_2759_, w_1923_, w_2692_);
and (w_0730_, w_1842_, w_1474_);
and (w_2755_, w_2069_, w_0517_);
and (w_1371_, w_3140_, w_1432_);
or (w_1754_, w_0714_, w_3378_);
or (w_3455_, w_1313_, w_3400_);
or (w_1470_, w_0499_, w_2151_);
or (out19[2], w_1242_, w_2740_);
not (w_1328_, w_2406_);
or (out11[1], w_1117_, w_3395_);
and (w_2266_, w_2966_, w_3217_);
not (w_3081_, w_1495_);
not (w_3266_, w_1293_);
or (w_3095_, w_1088_, w_2183_);
and (w_0024_, in3[1], w_0830_);
or (w_0845_, in11[6], w_1465_);
not (w_0934_, w_1253_);
and (w_3152_, in3[4], w_1363_);
or (w_1990_, w_0260_, w_2683_);
or (w_2333_, w_1348_, w_1524_);
or (w_2448_, w_2719_, w_2373_);
and (w_1026_, w_0790_, w_3330_);
or (w_3372_, w_0658_, w_0237_);
or (w_0755_, w_0607_, w_1804_);
not (w_3073_, in8[3]);
not (w_0136_, w_2050_);
or (w_1641_, w_0276_, w_2284_);
and (w_1156_, w_1028_, w_0163_);
or (w_1020_, w_0211_, w_0898_);
not (w_1715_, w_0973_);
not (w_0878_, w_1742_);
not (w_2517_, w_0671_);
or (w_0678_, in3[3], w_2892_);
or (w_2636_, w_0962_, w_1226_);
not (w_2181_, w_0965_);
or (w_1894_, w_3356_, w_3232_);
or (out23[3], w_1962_, w_1884_);
and (out13[4], w_1051_, w_2681_);
and (out24[7], w_2794_, w_1847_);
and (w_2108_, in14[0], w_2094_);
not (w_2463_, w_3014_);
and (w_2167_, out13[6], w_1808_);
and (w_3390_, in11[2], w_1703_);
and (w_0309_, w_1317_, w_2675_);
and (w_3096_, w_0608_, w_1826_);
and (w_0575_, w_2690_, w_0243_);
or (w_1706_, w_1744_, w_1499_);
or (w_1211_, w_3309_, w_0600_);
or (w_2018_, in15[2], w_2176_);
not (w_0686_, w_2865_);
or (w_2338_, w_1356_, w_2986_);
and (w_3197_, w_2175_, w_0693_);
and (w_2113_, in3[5], w_1531_);
or (w_2403_, in4[4], w_0765_);
and (w_1143_, w_0790_, w_3021_);
not (w_0704_, w_1244_);
or (w_2196_, w_1081_, w_0980_);
not (w_0200_, w_3328_);
or (w_0036_, w_2474_, w_1128_);
and (w_3352_, w_2162_, w_3344_);
not (w_1010_, in6[0]);
and (w_1663_, w_0915_, w_2925_);
or (w_0572_, w_2566_, w_1696_);
or (w_2904_, w_0907_, w_3030_);
and (w_0649_, w_2516_, w_3102_);
not (w_0861_, w_1626_);
not (w_3272_, w_0585_);
or (w_1162_, w_0599_, w_3228_);
or (w_0277_, w_1628_, w_2396_);
or (w_1448_, w_0694_, w_2182_);
not (w_0483_, w_2127_);
or (w_0995_, w_3007_, w_0238_);
and (w_2879_, w_0112_, w_0992_);
or (w_1234_, w_2223_, w_3255_);
and (w_0636_, w_3183_, w_3248_);
or (w_1504_, w_0730_, w_2660_);
or (w_0676_, w_1010_, w_2998_);
or (w_1937_, w_0291_, w_1685_);
or (w_1007_, w_1763_, w_3471_);
and (w_1711_, w_2888_, w_0957_);
or (w_1912_, w_1834_, w_2582_);
or (w_1353_, w_1474_, w_3175_);
and (w_1730_, w_2199_, w_1546_);
or (w_1480_, w_3205_, w_2382_);
and (w_0537_, w_0807_, w_1780_);
or (w_0050_, w_0317_, w_3113_);
or (w_1564_, w_3510_, w_1767_);
or (w_3526_, w_0952_, w_0182_);
and (w_3368_, in12[0], w_2745_);
not (w_0158_, w_2636_);
and (w_3346_, w_0005_, w_3086_);
and (w_1617_, w_0383_, w_0150_);
and (w_2975_, w_0488_, w_3249_);
and (w_2153_, w_2245_, w_2187_);
and (w_2730_, w_0233_, w_2823_);
and (w_2865_, in14[6], in13[6]);
or (w_0977_, w_2772_, w_0267_);
not (w_1900_, w_2990_);
or (w_1685_, w_2321_, w_0335_);
not (w_1577_, w_1807_);
and (w_1585_, w_1468_, w_0979_);
not (w_0394_, w_0356_);
and (w_1076_, w_2811_, w_0610_);
or (w_2990_, w_0669_, w_1987_);
not (w_0843_, w_1034_);
or (w_1229_, in13[0], w_0196_);
and (w_1296_, w_2095_, w_1135_);
or (w_3429_, w_0508_, w_1895_);
and (w_2139_, w_1294_, w_2904_);
and (w_2969_, w_1452_, w_3426_);
not (w_3173_, w_0192_);
and (out22[3], w_1184_, w_3245_);
or (w_1180_, w_1495_, w_2279_);
or (w_2508_, w_3405_, w_1383_);
not (w_0138_, in12[3]);
or (w_1202_, w_1286_, w_1799_);
and (w_2954_, w_2144_, w_2513_);
not (w_0119_, w_1427_);
not (w_0040_, w_3391_);
or (w_2613_, w_3345_, w_0242_);
or (w_1832_, in16[0], w_3079_);
and (w_1739_, w_0009_, w_2379_);
or (w_2626_, w_3153_, w_2705_);
and (w_3425_, w_2841_, w_2498_);
and (w_1819_, w_2019_, w_2153_);
and (w_0663_, w_1616_, w_1519_);
or (w_0305_, w_3179_, w_1924_);
or (w_1589_, w_2474_, w_1750_);
or (w_1028_, w_2955_, w_2320_);
or (w_2664_, w_2803_, w_3297_);
and (w_1927_, w_0658_, w_0237_);
or (out15[0], w_2572_, w_0100_);
or (w_1198_, w_1853_, w_1624_);
and (w_1872_, w_0277_, w_2812_);
and (w_1526_, w_0421_, w_3528_);
or (w_0919_, w_0730_, w_0638_);
and (w_2418_, w_1436_, w_1531_);
or (w_2084_, in7[5], w_1571_);
and (w_1155_, in14[6], w_3103_);
or (w_1032_, w_2175_, w_0418_);
not (w_3166_, w_2747_);
or (w_2109_, w_2961_, w_1192_);
or (w_1182_, w_1982_, w_1613_);
or (w_0681_, w_1095_, w_2073_);
and (w_0918_, w_0499_, w_2151_);
and (w_3052_, w_0941_, w_3371_);
and (w_1834_, w_1694_, w_1699_);
and (w_2938_, w_2658_, w_0658_);
and (w_0478_, w_0247_, w_3517_);
or (w_0951_, in14[0], w_2094_);
or (w_0179_, w_0793_, w_0279_);
or (w_2498_, w_2233_, w_0393_);
or (w_0842_, w_2414_, w_2869_);
or (w_2601_, in14[4], in13[4]);
or (w_1488_, in9[4], in10[0]);
and (w_2385_, w_2579_, w_3481_);
or (w_2840_, in16[7], in15[7]);
or (w_2987_, w_0796_, w_0856_);
and (w_0773_, w_0097_, w_1702_);
or (w_0406_, w_2417_, w_3461_);
not (w_3182_, w_0260_);
and (w_2388_, w_2670_, w_0911_);
or (w_1865_, w_1597_, w_1942_);
and (w_2161_, w_0363_, w_3138_);
and (w_1222_, w_1673_, w_2518_);
or (w_1909_, w_1870_, w_1642_);
and (w_1309_, w_2532_, w_1600_);
and (w_2933_, w_2249_, w_0083_);
not (w_1273_, w_2042_);
or (w_1333_, in9[5], in10[5]);
and (out21[3], w_1973_, w_3504_);
or (w_0130_, w_0808_, w_1920_);
and (w_2555_, in15[3], w_1618_);
or (w_0257_, w_0351_, w_1414_);
and (w_2767_, w_1742_, w_2784_);
or (w_0612_, w_3279_, w_3289_);
or (w_1722_, w_3484_, w_0435_);
or (w_3080_, w_0666_, w_2343_);
and (w_1948_, w_2995_, w_2331_);
and (w_2251_, w_2571_, w_0110_);
or (w_1702_, in3[5], w_2195_);
or (w_2422_, in14[2], in13[2]);
and (w_3412_, w_3469_, w_0691_);
or (w_2824_, w_1787_, w_0567_);
or (out16[5], w_0398_, w_2575_);
and (w_0854_, w_0132_, w_0451_);
or (w_2819_, w_0106_, w_3210_);
and (w_1110_, w_0836_, w_0286_);
and (w_2230_, w_2493_, w_0411_);
and (w_2963_, w_1716_, w_1171_);
or (w_1540_, w_0120_, w_0103_);
and (w_0434_, w_2253_, w_2454_);
or (w_1084_, w_1883_, w_2988_);
or (w_1800_, w_1144_, w_1475_);
and (w_1403_, w_2129_, w_0068_);
and (w_3456_, w_0187_, w_0251_);
or (w_0924_, w_2202_, w_0146_);
and (w_2502_, w_1590_, w_3237_);
not (w_1375_, w_0589_);
or (w_1388_, w_2967_, w_3502_);
and (w_2910_, in13[5], w_3359_);
or (w_2405_, w_2931_, w_2810_);
or (w_3055_, w_0548_, w_1116_);
or (w_3044_, in8[3], w_1397_);
or (w_0611_, w_2421_, w_3266_);
and (w_0367_, w_0599_, w_1588_);
or (w_3083_, in6[0], w_3134_);
and (out17[7], w_2371_, w_0873_);
and (w_1144_, w_0421_, w_2338_);
and (w_1880_, w_3352_, w_0271_);
or (w_2170_, w_1932_, w_3053_);
or (w_1886_, w_0175_, w_1252_);
and (w_2489_, w_2451_, w_0972_);
and (w_0126_, w_0064_, w_2356_);
or (w_2215_, w_1607_, out13[2]);
and (w_2033_, w_2961_, w_1675_);
or (w_1859_, w_2579_, w_3481_);
or (w_0472_, w_2959_, w_0281_);
and (out14[5], w_1757_, w_3373_);
or (w_3187_, w_1466_, w_1030_);
or (w_0820_, w_1460_, w_1523_);
and (w_0146_, w_1527_, w_1481_);
and (w_0180_, w_2163_, w_3468_);
not (w_3301_, w_2113_);
not (w_0960_, in6[5]);
or (w_2024_, in4[4], w_1611_);
or (w_2288_, w_2828_, w_1138_);
and (out7[3], w_2594_, w_2573_);
and (w_0369_, w_3352_, w_3051_);
or (w_0003_, w_0814_, w_2430_);
or (w_1224_, w_2563_, w_3021_);
and (w_2914_, w_3154_, w_2443_);
and (out2[1], w_2636_, w_2561_);
not (w_3405_, w_1429_);
or (w_3314_, w_2227_, w_0422_);
or (w_1276_, w_2228_, w_0828_);
and (w_0808_, w_2936_, w_2333_);
or (w_3119_, in13[7], w_3038_);
and (w_1964_, w_0521_, w_3109_);
and (w_1301_, in15[7], w_2764_);
or (w_0137_, w_0616_, w_2634_);
or (w_0917_, w_2959_, w_2009_);
not (w_0789_, w_2167_);
or (w_1683_, w_2917_, w_1342_);
or (w_0193_, in16[5], w_0090_);
not (w_1235_, w_1224_);
or (out5[3], w_3313_, w_1222_);
and (w_3065_, w_3261_, w_1079_);
not (w_1137_, w_1692_);
and (w_3170_, w_1714_, w_0747_);
and (w_0428_, w_3405_, w_1150_);
or (w_3325_, w_0963_, w_1977_);
or (w_1527_, w_3484_, w_1113_);
not (w_1099_, w_1462_);
and (w_0323_, w_1398_, w_0575_);
or (w_1129_, in12[7], w_2651_);
or (w_2594_, w_3108_, w_3284_);
or (w_1324_, w_1066_, w_0352_);
or (w_0159_, w_2976_, w_0360_);
or (w_3335_, w_0617_, w_3459_);
and (w_2934_, w_1660_, w_1347_);
or (w_2695_, w_2135_, w_1137_);
or (w_0354_, w_2415_, w_2068_);
or (w_2886_, w_1680_, w_1181_);
and (w_2639_, w_1859_, w_0257_);
not (w_0584_, w_2038_);
or (w_2925_, w_0687_, w_1092_);
or (w_0445_, w_2390_, w_1072_);
or (out15[3], w_1838_, w_0288_);
or (w_1056_, w_3253_, w_0180_);
and (w_3435_, w_1208_, w_1938_);
and (w_0914_, w_0034_, w_1174_);
not (w_0155_, w_0411_);
and (w_1104_, w_0421_, w_0456_);
and (w_1150_, w_1153_, w_0145_);
or (w_2101_, w_2650_, w_2390_);
and (w_2817_, w_1843_, w_2623_);
not (w_0427_, w_0689_);
and (w_0607_, w_3328_, w_3183_);
and (w_2762_, w_2447_, w_0716_);
and (w_3209_, w_3186_, w_0647_);
or (w_2532_, w_1041_, w_1002_);
and (w_0523_, w_1084_, w_0776_);
and (w_0877_, w_0666_, w_1030_);
and (w_0298_, w_0453_, w_2011_);
or (w_1409_, w_2959_, w_0407_);
and (w_1758_, in8[0], w_1238_);
or (w_1280_, w_0927_, w_2476_);
or (w_1125_, w_0990_, w_0773_);
or (w_2187_, w_1639_, w_1338_);
not (w_2598_, w_3412_);
and (w_0769_, w_2635_, w_0147_);
or (w_0568_, w_0458_, w_2829_);
and (w_2445_, w_2014_, w_2993_);
not (w_1390_, w_1725_);
not (w_3048_, in7[5]);
or (w_0925_, w_0390_, w_1148_);
not (w_0703_, out16[1]);
not (w_0644_, w_0143_);
or (w_0065_, w_0690_, w_0637_);
or (w_0124_, w_2795_, w_3464_);
and (w_2541_, w_2370_, w_1307_);
and (w_2546_, in14[1], in13[1]);
and (out10[2], w_1416_, w_3299_);
or (w_1416_, w_1736_, w_1008_);
and (w_3480_, w_0550_, w_2381_);
or (w_3489_, w_1965_, w_2329_);
and (w_0544_, w_3111_, w_3120_);
or (w_2521_, in7[0], w_2023_);
or (w_0173_, w_0700_, w_1913_);
and (w_2711_, w_1429_, w_1466_);
or (w_2371_, w_1663_, w_1881_);
and (w_3190_, w_2859_, w_1543_);
not (w_0127_, w_1214_);
and (w_1972_, w_3153_, w_2705_);
or (w_0930_, w_0096_, w_1012_);
or (w_3241_, w_1455_, w_2543_);
or (w_1915_, in1[1], in2[2]);
or (w_2379_, w_1654_, w_2006_);
and (out15[6], w_1233_, w_1496_);
or (w_0234_, w_2487_, w_0724_);
and (w_2377_, w_3375_, w_3403_);
and (w_2252_, w_0892_, w_0651_);
or (w_2332_, in1[3], in2[3]);
not (w_1605_, in8[1]);
or (w_2974_, w_0942_, w_3501_);
or (w_3029_, w_0341_, w_3252_);
or (w_0097_, w_0215_, w_2434_);
and (w_1053_, w_1033_, w_1551_);
not (w_2750_, w_1373_);
and (w_0260_, w_0214_, w_2637_);
or (w_2070_, w_1519_, w_2057_);
and (w_1376_, w_2467_, w_0955_);
and (w_2098_, w_2942_, w_1060_);
and (w_0654_, w_0781_, w_3528_);
or (out11[5], w_0080_, w_3087_);
or (w_2580_, w_2934_, w_0771_);
and (w_3228_, w_1877_, w_0372_);
and (w_2618_, w_0823_, w_2446_);
and (w_0096_, w_2494_, w_1899_);
or (w_1707_, w_0188_, w_1352_);
and (out4[3], w_2491_, w_0406_);
or (w_2687_, w_0639_, w_0505_);
or (w_2655_, w_0942_, w_0060_);
and (w_2778_, w_1815_, w_0939_);
and (w_2869_, w_2169_, w_2071_);
not (w_2000_, in1[2]);
not (w_2658_, w_3172_);
and (w_0268_, w_1057_, w_3116_);
not (w_3199_, in15[4]);
and (w_2277_, w_2717_, w_3059_);
or (w_1316_, w_2952_, w_0821_);
or (w_0848_, w_3329_, w_3191_);
or (w_0884_, w_0993_, w_1606_);
or (w_2124_, w_2207_, w_0333_);
or (w_1418_, w_0657_, w_2791_);
or (w_2162_, w_0603_, w_0874_);
and (w_1261_, w_1488_, w_0081_);
not (w_0052_, w_0332_);
and (w_1354_, w_1698_, w_0511_);
and (w_3528_, w_1690_, w_3301_);
and (w_2846_, w_0137_, w_0507_);
and (w_3442_, w_2888_, w_2062_);
or (w_0511_, w_2613_, w_0677_);
and (w_2453_, w_3469_, w_1494_);
and (out15[4], w_0167_, w_2997_);
not (w_0959_, w_3071_);
or (w_3229_, w_2665_, w_1059_);
and (w_0765_, w_1085_, w_2273_);
and (w_0520_, w_2803_, w_3297_);
and (w_0879_, w_2673_, w_1370_);
or (w_2993_, w_0133_, w_1385_);
and (w_2298_, w_1190_, w_2126_);
or (w_0328_, w_1485_, w_2496_);
or (w_2874_, w_2153_, w_3105_);
or (w_3230_, in11[1], w_0965_);
not (w_2896_, w_1060_);
or (w_3468_, w_1558_, w_2246_);
or (w_3391_, w_1227_, w_2208_);
not (w_2796_, in13[4]);
and (w_0249_, w_2955_, w_0322_);
or (w_1021_, w_1429_, w_3510_);
and (w_1753_, w_3060_, w_0434_);
not (w_1245_, w_3466_);
and (w_1254_, w_3262_, w_2168_);
and (w_2490_, w_2792_, w_3476_);
or (w_3353_, w_0441_, w_0361_);
not (w_0542_, w_1606_);
and (w_0598_, w_1491_, w_3033_);
or (w_3126_, w_2121_, w_3516_);
not (w_2413_, in15[5]);
or (w_1188_, w_0599_, w_1588_);
and (w_1652_, w_1401_, w_2398_);
and (w_3322_, w_0708_, w_2947_);
or (w_1591_, w_0688_, w_2356_);
not (w_1361_, in1[4]);
and (w_3045_, w_2967_, w_3502_);
and (w_2588_, in11[7], w_0884_);
or (w_2737_, out13[6], w_1808_);
and (w_0630_, w_1315_, in13[5]);
or (w_0442_, w_1025_, w_3343_);
and (w_1762_, w_2319_, w_2859_);
and (out10[4], w_2786_, w_1101_);
not (w_0910_, w_0069_);
and (out9[4], w_2464_, w_0494_);
or (w_2916_, w_3278_, w_2497_);
and (w_0390_, w_2563_, w_1616_);
not (w_2157_, w_0347_);
not (w_2895_, w_0942_);
not (w_1877_, w_1519_);
and (w_1622_, in11[5], w_3479_);
or (out20[0], w_1550_, w_3490_);
and (w_0088_, w_1861_, w_1837_);
and (w_3090_, w_0676_, w_3083_);
and (w_3196_, w_2566_, w_1696_);
or (w_1086_, in7[1], w_2200_);
and (out6[1], w_1616_, w_3218_);
and (w_1561_, w_2312_, w_0071_);
or (w_2669_, w_0282_, w_0858_);
or (out4[5], w_3065_, w_0077_);
and (w_3366_, w_0521_, w_0193_);
or (w_2739_, w_0122_, w_3258_);
and (w_0484_, w_0123_, w_0270_);
or (w_1898_, w_1862_, w_0030_);
and (w_0557_, w_3454_, w_0640_);
not (w_1106_, w_2897_);
or (w_2350_, out14[5], w_1761_);
and (w_2200_, w_2147_, w_2697_);
and (w_0062_, w_1651_, w_1877_);
and (w_0244_, w_3241_, w_1540_);
or (w_1679_, w_0520_, w_2558_);
or (w_2056_, w_0562_, w_1260_);
or (w_0795_, w_0387_, w_1873_);
and (w_1077_, w_0237_, w_3435_);
or (out18[1], w_3034_, w_0237_);
not (w_1511_, w_0607_);
not (w_1563_, w_1094_);
not (w_3261_, w_0205_);
or (w_2147_, w_0676_, w_1709_);
not (w_0700_, w_0241_);
and (w_1727_, w_0849_, w_3143_);
or (w_1377_, w_2580_, w_3263_);
and (w_0226_, w_3367_, w_2047_);
and (w_1635_, w_2206_, w_0416_);
or (w_0946_, w_2817_, w_1247_);
or (w_2245_, w_0544_, w_1816_);
and (w_3451_, w_1892_, w_0350_);
not (w_2749_, w_3196_);
or (w_2530_, w_3297_, w_0760_);
or (w_2793_, w_0268_, w_3180_);
or (w_2701_, w_0089_, w_2181_);
and (w_1181_, w_0652_, w_2500_);
or (out18[6], w_1535_, w_3060_);
or (w_1543_, w_2285_, w_3099_);
and (w_2173_, w_3114_, w_2056_);
or (w_0812_, w_2501_, w_3451_);
or (w_1716_, w_0099_, w_1449_);
and (w_0983_, w_0365_, w_2275_);
and (w_1867_, w_0800_, w_3351_);
and (w_3007_, w_0217_, w_0244_);
not (w_2428_, w_0879_);
and (w_2473_, w_0666_, w_0221_);
or (w_2890_, in7[1], w_3163_);
or (w_0005_, w_3267_, w_3084_);
or (w_2441_, w_0893_, w_0021_);
and (w_1126_, w_1491_, w_3522_);
or (w_1011_, w_3218_, w_0781_);
or (w_1733_, w_1770_, w_2044_);
and (w_0952_, in15[5], w_2100_);
and (w_3415_, w_0568_, w_1165_);
or (w_1950_, w_0142_, w_0880_);
and (w_1884_, w_1308_, w_2119_);
and (w_2595_, w_0035_, w_2356_);
and (w_3192_, in14[2], w_3420_);
or (w_1933_, w_3368_, w_2224_);
not (w_0026_, w_2018_);
and (w_2430_, w_0112_, w_0510_);
and (w_0891_, w_3267_, w_1174_);
or (w_1055_, w_2815_, w_2965_);
or (w_0881_, w_2193_, w_2053_);
or (w_2436_, w_0491_, w_0373_);
or (w_3396_, w_0786_, w_1375_);
or (w_1878_, w_3225_, w_1107_);
not (w_3279_, w_1274_);
and (w_0740_, w_1284_, w_3098_);
and (w_1669_, w_3487_, w_1126_);
and (w_3496_, in1[4], in2[5]);
and (w_2482_, w_0395_, w_0203_);
and (w_2006_, w_2923_, w_1258_);
and (w_2064_, w_3109_, w_2103_);
or (w_3344_, w_0614_, w_0292_);
and (w_0319_, w_2959_, w_1401_);
not (w_0056_, w_3263_);
not (w_3463_, w_3077_);
or (w_2923_, w_1901_, w_3196_);
or (w_0899_, w_2755_, w_1793_);
or (w_0803_, w_1992_, w_3407_);
or (w_2126_, w_2843_, w_0859_);
or (w_1544_, w_1043_, w_0108_);
or (w_1764_, w_0480_, w_2774_);
or (w_0488_, w_0582_, w_1197_);
or (w_2278_, w_2175_, w_0217_);
or (w_0389_, w_0290_, w_2355_);
or (w_2020_, w_2383_, w_3181_);
not (w_2105_, w_2508_);
and (w_2538_, w_3297_, w_1220_);
and (w_0941_, w_2206_, w_2178_);
and (out10[1], w_1766_, w_0925_);
and (w_3323_, w_3200_, w_3150_);
and (w_0175_, in3[3], w_0266_);
or (w_2396_, w_1893_, w_0819_);
or (w_1398_, w_2851_, w_1744_);
and (w_2753_, w_1313_, w_3400_);
or (w_0844_, w_1206_, w_2048_);
or (w_0939_, w_1127_, out13[1]);
or (w_0141_, w_2629_, w_2267_);
and (w_1959_, w_1992_, w_3407_);
or (w_1172_, in3[4], w_1363_);
or (w_1124_, w_0061_, w_3238_);
or (w_2419_, w_2499_, w_1733_);
and (w_2699_, w_3507_, w_1852_);
and (w_2863_, w_1764_, w_1687_);
or (w_3121_, in15[5], in16[5]);
or (w_1700_, w_3157_, w_2287_);
or (w_0163_, w_3049_, w_0874_);
not (w_3285_, w_2991_);
and (out6[3], w_2563_, w_3105_);
or (w_3105_, w_2903_, w_2884_);
and (w_0800_, w_2990_, w_2237_);
and (w_0661_, w_3473_, w_1833_);
or (w_0631_, w_2065_, w_2850_);
and (out9[2], w_1268_, w_0047_);
or (w_2265_, w_0214_, w_2637_);
not (w_3518_, w_3522_);
and (w_1523_, w_3288_, w_1762_);
not (w_2912_, w_2842_);
not (w_2516_, w_1771_);
or (w_1742_, w_2292_, w_2979_);
and (w_3210_, w_1435_, w_3133_);
or (w_3145_, w_0317_, w_2798_);
or (w_1776_, w_3501_, w_0064_);
and (w_3490_, w_1466_, w_1277_);
or (w_2012_, w_1493_, w_0623_);
not (w_1256_, w_1913_);
and (w_2900_, w_0790_, w_0599_);
and (w_0958_, w_1141_, w_3501_);
or (w_3032_, w_0469_, w_1947_);
and (w_0660_, w_0480_, w_2774_);
and (w_0690_, w_0500_, w_1973_);
and (w_1091_, in14[4], w_3466_);
not (w_1719_, w_0034_);
and (w_1072_, w_0546_, w_1889_);
and (w_1330_, w_1127_, out13[1]);
not (w_1436_, w_3034_);
or (w_0954_, w_0942_, w_0848_);
or (w_0811_, w_0661_, w_1310_);
or (w_3311_, in11[3], w_0643_);
and (w_1971_, in7[4], w_0833_);
and (w_0424_, w_0609_, w_0051_);
or (w_0519_, w_0138_, w_2750_);
and (w_0763_, w_3187_, w_2225_);
or (w_2232_, w_0161_, w_0504_);
or (w_2549_, w_2362_, w_0062_);
and (w_0123_, w_0272_, w_0094_);
or (w_1196_, w_0790_, w_3385_);
or (w_0620_, w_1830_, w_2603_);
or (w_2244_, w_1325_, w_2131_);
and (w_1019_, w_2814_, w_2122_);
and (w_2892_, w_1090_, w_0050_);
or (w_0882_, w_2108_, w_2201_);
or (w_0945_, w_0376_, w_0731_);
and (w_2057_, w_1742_, w_1846_);
not (w_1556_, w_2460_);
and (w_0720_, w_2722_, w_1872_);
or (w_1164_, w_1971_, w_2878_);
not (w_0626_, w_2174_);
or (w_2535_, w_2479_, w_1195_);
and (w_1606_, in9[7], in10[3]);
and (w_0455_, w_1768_, w_0151_);
or (w_3089_, w_3336_, w_2804_);
or (w_1334_, in11[7], w_1822_);
and (w_2671_, w_0255_, w_1372_);
and (w_1699_, w_1995_, w_2655_);
and (w_0220_, in6[5], in5[4]);
and (w_2792_, w_1538_, w_1360_);
or (w_2607_, w_3510_, out13[0]);
and (w_1413_, w_1401_, w_0844_);
and (w_2145_, w_1171_, w_2158_);
or (w_1714_, w_0912_, w_1272_);
and (w_3497_, w_0116_, w_1829_);
or (w_3138_, w_2185_, w_1030_);
or (w_0112_, w_2096_, w_0381_);
or (w_1360_, w_1139_, w_3047_);
or (w_3072_, in12[3], w_1373_);
and (w_0745_, w_3034_, w_3293_);
or (out23[2], w_2822_, w_1559_);
and (w_0357_, w_0121_, w_0529_);
or (w_3017_, w_3510_, w_1495_);
or (w_1766_, w_0079_, w_2088_);
or (w_3116_, w_0722_, w_3270_);
and (w_0402_, out9[0], w_2968_);
or (w_1588_, w_0711_, w_0498_);
and (w_1535_, w_3383_, w_2160_);
and (w_0938_, w_1325_, w_2898_);
not (w_1329_, w_0064_);
or (w_1167_, in11[7], w_0884_);
and (w_3103_, w_1050_, w_2562_);
or (w_0894_, w_0152_, w_1972_);
and (w_1807_, w_0466_, w_1303_);
or (w_2550_, w_0665_, w_1281_);
or (w_3185_, in16[3], w_0818_);
and (w_3123_, w_1814_, out16[2]);
not (w_1713_, w_3052_);
not (w_0002_, w_2570_);
and (w_2785_, w_3156_, w_2628_);
and (w_2769_, w_3023_, w_2328_);
and (w_2325_, w_1368_, w_1321_);
not (w_2596_, w_1631_);
or (w_0999_, w_2052_, w_1450_);
or (w_1300_, w_1390_, w_2865_);
and (w_1358_, w_3415_, w_0587_);
not (w_2630_, w_1265_);
or (w_2014_, w_2059_, w_1797_);
and (w_2361_, w_2980_, w_0447_);
and (w_2971_, w_0471_, w_2052_);
and (w_2845_, w_0961_, w_0358_);
not (w_2809_, w_1763_);
and (w_3458_, w_2009_, w_3269_);
or (w_2968_, w_0986_, w_1314_);
or (w_1984_, w_1340_, w_0670_);
or (w_0429_, w_3243_, w_1708_);
or (w_0012_, w_2172_, w_2897_);
and (w_1978_, in13[0], w_0196_);
and (out21[6], w_1826_, w_2395_);
or (w_3172_, w_2269_, w_3525_);
not (w_0134_, w_0838_);
not (w_2302_, in10[5]);
or (w_2380_, w_3229_, w_2357_);
not (w_2299_, w_1699_);
and (out17[4], w_0034_, w_0859_);
and (out17[2], w_0671_, w_3183_);
and (w_2534_, w_0351_, w_1414_);
and (w_2235_, in6[0], w_3134_);
not (w_1485_, w_2813_);
and (w_1130_, w_2629_, w_2267_);
not (w_1355_, w_0730_);
and (w_2893_, w_2402_, w_1704_);
or (w_0988_, w_1719_, w_1529_);
not (w_3041_, in14[6]);
and (w_1611_, w_2124_, w_0474_);
and (w_2205_, w_0960_, w_0497_);
or (w_0911_, w_0045_, w_2296_);
and (w_2263_, w_0023_, w_0038_);
not (w_0490_, w_1407_);
and (w_3134_, w_3139_, w_0475_);
not (w_2198_, out9[0]);
or (w_1184_, w_2289_, w_2714_);
or (w_1637_, w_2609_, w_0934_);
not (w_1534_, w_3404_);
or (w_0121_, w_2630_, w_0768_);
and (out14[1], w_0589_, w_2920_);
or (w_3443_, w_2567_, w_0810_);
or (w_3434_, w_1483_, w_1718_);
or (w_0827_, w_2061_, w_1302_);
and (w_1810_, w_1440_, w_2663_);
not (w_0451_, w_3351_);
and (w_1238_, w_0438_, w_0668_);
and (w_0896_, w_1768_, w_0303_);
or (w_0841_, w_3445_, w_3094_);
and (w_0131_, w_1139_, w_3047_);
or (w_2760_, w_0151_, w_2299_);
or (w_1516_, w_0555_, w_3011_);
or (w_1121_, w_0615_, w_3508_);
or (w_1449_, w_1107_, w_0484_);
and (w_3071_, w_3182_, w_2265_);
and (w_1840_, w_0233_, w_0140_);
not (w_2449_, out14[7]);
not (w_0133_, w_2223_);
or (out5[4], w_2711_, w_0428_);
and (w_2402_, in7[0], w_3090_);
and (w_1127_, w_0666_, w_0271_);
or (w_2319_, w_2086_, w_2827_);
and (w_2628_, w_0888_, w_2964_);
or (w_1920_, w_1437_, w_0983_);
and (w_1338_, w_0286_, w_0648_);
or (w_1147_, w_0048_, w_1261_);
or (w_3148_, w_2009_, w_2266_);
not (w_1288_, w_1840_);
or (w_2416_, w_3199_, w_1111_);
or (out8[1], w_0745_, w_3193_);
or (w_3260_, in6[1], w_0872_);
or (w_0310_, in1[2], in2[3]);
not (w_1802_, w_1314_);
or (w_1050_, w_3318_, w_1722_);
or (w_3294_, w_2064_, w_3352_);
or (w_1339_, w_2173_, w_3068_);
or (w_1492_, w_0253_, w_3024_);
or (w_2192_, w_3330_, w_2669_);
and (w_0344_, w_1909_, w_3176_);
or (w_0094_, w_2146_, w_0306_);
not (w_1858_, w_1931_);
and (w_2575_, w_1877_, w_3330_);
and (w_3483_, w_0257_, w_2239_);
or (w_0029_, w_3014_, w_1331_);
or (w_0897_, in1[0], in2[0]);
or (w_3375_, w_0514_, w_0483_);
not (w_2097_, w_2745_);
or (w_3104_, in8[4], w_2751_);
and (w_0192_, w_1498_, w_3075_);
or (w_0364_, in9[0], in10[0]);
or (w_2500_, in7[4], w_0833_);
and (w_2758_, w_0034_, w_2086_);
and (w_2315_, w_1429_, w_0599_);
or (w_1336_, w_0059_, w_2733_);
and (out21[1], w_2293_, w_3273_);
and (w_1731_, w_3510_, w_1401_);
not (w_2775_, w_0746_);
not (w_2657_, out16[7]);
and (w_2850_, w_0562_, w_1260_);
and (w_0597_, w_1044_, w_1037_);
or (w_2440_, w_1771_, w_0799_);
not (w_3097_, w_1476_);
and (w_2552_, in3[1], w_2666_);
or (out14[7], w_0762_, w_3274_);
and (w_0240_, w_1190_, w_2908_);
and (w_2600_, w_0229_, w_1120_);
and (w_2578_, in9[3], in10[3]);
and (w_0223_, w_0841_, w_1133_);
or (w_3254_, in7[2], w_1311_);
and (w_2909_, w_0388_, w_1004_);
and (w_2853_, w_0271_, w_3297_);
and (w_2915_, w_3229_, w_2357_);
or (w_0303_, w_2827_, w_1625_);
and (w_1192_, w_2908_, w_1575_);
and (w_0282_, w_3283_, w_2946_);
not (w_0880_, w_1672_);
and (w_2646_, w_0804_, w_0658_);
or (w_1520_, w_3149_, w_2220_);
and (w_2352_, w_3114_, w_2899_);
or (w_0696_, w_2163_, w_3468_);
and (out16[1], w_1875_, w_3372_);
or (w_2935_, w_1720_, w_1941_);
not (w_0864_, w_3379_);
or (w_0431_, w_3023_, w_2328_);
and (w_3330_, w_1062_, w_1713_);
or (w_1583_, w_1562_, w_0936_);
or (w_2229_, w_0119_, w_0220_);
and (w_3498_, in11[6], w_1237_);
and (w_2612_, w_1661_, w_2462_);
not (w_3478_, w_2776_);
and (w_0106_, in1[2], in2[2]);
or (w_0707_, w_1668_, w_2785_);
or (w_0733_, w_0329_, w_0154_);
and (w_1369_, w_2013_, w_3029_);
and (w_1787_, in5[2], w_2063_);
and (w_2093_, w_1538_, w_0678_);
and (w_2733_, w_3470_, w_1251_);
and (w_2725_, w_0519_, w_3200_);
or (w_3046_, w_2837_, w_1841_);
or (w_3033_, w_2456_, w_3025_);
or (w_3439_, w_1574_, w_3045_);
and (w_2001_, w_1043_, w_0108_);
and (w_0258_, w_1015_, w_1339_);
or (w_1134_, w_2307_, w_1351_);
and (w_0346_, in13[3], w_3323_);
or (w_2557_, w_2832_, w_3342_);
and (w_0152_, in16[3], w_0818_);
and (w_3411_, w_0416_, w_1895_);
and (w_1696_, w_0212_, w_1162_);
or (w_2722_, w_3331_, w_0524_);
and (w_1601_, w_0966_, w_3260_);
or (w_3220_, in14[1], in13[1]);
and (w_0460_, w_0840_, w_2424_);
or (w_2898_, w_0943_, w_1519_);
not (w_0605_, w_1132_);
or (w_1173_, w_0622_, w_0875_);
or (w_0990_, w_1595_, w_0720_);
not (w_3002_, w_2487_);
not (w_3076_, w_0768_);
and (w_0007_, in14[5], w_2777_);
or (w_0521_, w_1443_, w_0371_);
and (out4[0], w_1547_, w_1998_);
and (w_1022_, w_3043_, w_0213_);
or (w_3306_, w_0685_, w_0883_);
and (w_3413_, w_3108_, w_1677_);
or (w_2412_, w_2595_, w_2620_);
or (w_1725_, in14[6], in13[6]);
not (w_1102_, w_1869_);
or (w_2485_, w_0183_, w_1684_);
and (w_3281_, w_2810_, w_0624_);
and (w_1839_, w_0326_, w_1094_);
or (w_3231_, w_1301_, w_2537_);
not (w_2225_, w_0171_);
and (w_0832_, w_2213_, w_1248_);
and (w_2094_, w_1813_, w_1229_);
and (w_0558_, w_3073_, w_1023_);
and (w_3505_, in7[1], w_2200_);
or (w_2706_, w_3124_, w_0601_);
not (w_2529_, w_1627_);
not (w_1612_, w_3358_);
not (w_0048_, in11[4]);
not (w_1846_, w_2856_);
or (w_0207_, w_1964_, w_1364_);
or (w_2007_, w_2618_, w_0121_);
or (w_1487_, w_1617_, w_2915_);
and (w_2456_, w_1882_, w_1284_);
or (w_2406_, in11[4], w_3158_);
or (w_3461_, w_3453_, w_0767_);
or (w_0816_, in4[2], w_1930_);
not (w_1789_, w_3396_);
not (w_1216_, w_0914_);
and (w_3432_, w_2809_, w_1741_);
and (w_1793_, w_1991_, w_2255_);
and (w_0722_, w_0420_, w_1196_);
and (w_0407_, w_2807_, w_2747_);
or (w_2806_, w_2377_, w_2984_);
not (w_3360_, w_1809_);
not (w_1096_, w_2914_);
or (w_3290_, w_2509_, w_1905_);
and (w_1981_, in12[3], w_1373_);
and (w_1306_, w_3356_, w_3232_);
not (w_0974_, w_0202_);
or (w_2523_, w_1792_, w_0571_);
or (out3[3], w_1104_, w_1903_);
and (w_2179_, out14[2], w_1949_);
and (w_3258_, w_2944_, w_0827_);
and (out7[4], w_3314_, w_0812_);
or (w_3139_, w_2685_, w_1096_);
or (w_2218_, w_2533_, w_1478_);
or (w_3003_, w_1507_, w_0169_);
or (w_0213_, w_2852_, w_2412_);
and (w_0781_, w_2157_, w_0723_);
or (w_0829_, w_2566_, w_0859_);
or (w_0438_, w_3264_, w_1557_);
or (w_1345_, w_1616_, w_1519_);
or (w_1835_, w_2555_, w_1921_);
or (w_2953_, w_0137_, w_0507_);
or (w_0114_, w_2277_, w_1688_);
or (w_1892_, w_1719_, w_2820_);
and (out24[3], w_3365_, w_0719_);
not (w_3293_, w_3497_);
and (w_0480_, w_3234_, w_1243_);
or (w_3381_, w_1145_, w_1726_);
and (w_0090_, w_2781_, w_1943_);
and (w_2435_, w_1737_, w_3105_);
or (w_3403_, w_1813_, w_3488_);
not (w_2317_, w_2212_);
or (w_0218_, w_1616_, w_2545_);
and (w_1323_, w_3353_, w_0613_);
or (w_2045_, w_1280_, w_2410_);
and (w_3513_, in1[1], in2[2]);
or (w_0634_, w_2588_, w_1161_);
not (w_2300_, w_1581_);
or (w_2185_, w_0216_, w_0159_);
or (out23[6], w_0591_, w_0424_);
and (w_2082_, w_1471_, w_0561_);
not (w_3339_, w_3388_);
not (w_2519_, w_1152_);
and (w_3135_, w_0688_, w_2518_);
not (w_2553_, w_3410_);
and (w_2172_, w_3019_, w_2568_);
and (w_1991_, w_0652_, w_1640_);
not (w_1783_, w_2786_);
and (out17[0], w_0271_, w_2803_);
or (w_2814_, w_3498_, w_1669_);
and (w_2283_, in7[3], w_3257_);
or (w_3363_, w_0960_, w_0497_);
and (w_3426_, w_3315_, w_2349_);
or (w_0529_, w_1940_, w_2802_);
or (w_0153_, w_0301_, w_0437_);
or (w_3129_, w_0924_, w_1530_);
or (out8[0], w_2473_, w_0541_);
or (w_2906_, w_1720_, w_1925_);
and (w_3492_, w_1939_, w_1638_);
and (w_1967_, in11[4], w_3158_);
and (w_1750_, w_1381_, w_1216_);
and (w_2841_, w_0008_, w_2507_);
or (w_3521_, w_0249_, w_1515_);
not (w_3040_, w_1737_);
not (w_1777_, w_3138_);
not (w_0363_, w_1194_);
and (w_1067_, w_0420_, w_1057_);
not (w_0593_, w_3103_);
not (w_1383_, w_3060_);
and (w_0847_, w_2339_, w_0779_);
or (w_0043_, in14[2], w_3420_);
and (w_0157_, in16[7], in15[7]);
or (w_0892_, w_0543_, w_0230_);
or (w_2103_, w_3444_, w_3366_);
not (w_2998_, w_3134_);
and (w_1259_, w_3278_, w_2497_);
not (w_2714_, w_1990_);
not (w_2512_, in7[4]);
not (w_3326_, w_3121_);
or (w_0091_, w_2635_, w_0147_);
or (w_2743_, out15[0], w_2803_);
or (w_0471_, w_2957_, w_2418_);
and (w_0594_, w_2773_, w_2838_);
or (w_3188_, w_0329_, w_0642_);
and (w_0316_, w_1535_, w_3081_);
and (w_1970_, w_0421_, w_0631_);
and (w_1500_, w_2820_, w_0217_);
and (w_1619_, w_0162_, w_0389_);
or (w_2673_, w_1945_, w_1534_);
and (w_2901_, w_1058_, w_1778_);
and (w_2514_, in16[7], w_1462_);
and (out2[3], w_1801_, w_1225_);
and (w_2004_, w_1850_, w_2217_);
and (w_0064_, w_1377_, w_2698_);
or (w_1058_, w_3470_, w_1251_);
and (w_1720_, w_0181_, w_1457_);
and (w_0680_, w_2895_, w_0662_);
and (w_0871_, w_2827_, w_1625_);
and (w_1887_, w_0804_, w_3352_);
and (w_2271_, w_0501_, w_1895_);
or (w_1412_, w_1674_, w_0528_);
not (w_0463_, out14[3]);
or (w_0031_, w_3423_, w_1784_);
not (w_0462_, w_2625_);
and (w_1965_, w_0326_, w_2241_);
not (w_1266_, w_0504_);
and (w_0177_, out13[7], w_0929_);
and (w_2839_, w_0599_, w_1519_);
and (w_2092_, w_2518_, w_2009_);
not (w_0662_, w_1549_);
and (w_0922_, w_2038_, w_2827_);
or (w_3410_, w_0200_, w_2941_);
and (w_0017_, w_2459_, w_2565_);
and (w_3099_, w_2319_, w_0025_);
and (w_1097_, in15[5], in16[5]);
and (w_1350_, w_0482_, w_1898_);
not (w_2787_, w_3012_);
and (w_2060_, in16[4], w_3132_);
or (w_0243_, in4[2], w_2863_);
or (w_2130_, w_1194_, w_1777_);
or (w_2554_, w_3126_, w_0896_);
and (w_0895_, in4[3], w_1042_);
or (w_2838_, in13[6], w_2556_);
and (w_2528_, w_3375_, w_0549_);
or (w_1632_, w_3172_, w_3386_);
or (w_2622_, w_0852_, w_1460_);
not (w_0586_, w_2555_);
or (w_2583_, w_1854_, w_2569_);
and (w_0893_, in3[2], w_3280_);
or (w_2624_, w_2121_, w_3480_);
and (w_0486_, w_1348_, w_1524_);
and (w_2166_, w_3475_, w_1169_);
and (w_1308_, w_3510_, w_1519_);
not (w_1815_, w_1330_);
and (w_0535_, w_2422_, w_2186_);
or (w_1284_, w_2927_, w_0017_);
and (w_1936_, w_0550_, w_0999_);
not (w_0869_, w_1186_);
and (w_0975_, w_1544_, w_1276_);
or (w_1914_, w_2448_, w_2431_);
or (w_2746_, in11[4], w_1287_);
and (w_1694_, w_3126_, w_0896_);
and (w_0191_, w_0200_, w_2704_);
and (w_1454_, w_1175_, w_1017_);
and (w_1752_, w_2616_, w_2978_);
or (w_0420_, w_1673_, w_0712_);
or (w_0378_, in1[3], in2[4]);
or (out23[4], w_0414_, w_0540_);
and (w_0556_, w_0601_, w_0237_);
and (w_0739_, w_0908_, w_1532_);
or (w_0194_, w_3093_, w_0204_);
not (w_1357_, w_3359_);
or (w_2342_, w_1346_, w_1136_);
or (w_2679_, in4[5], w_1922_);
or (w_0652_, w_2512_, w_0445_);
or (w_1955_, w_3310_, w_2624_);
and (w_0468_, w_2523_, w_2031_);
or (w_1966_, w_2671_, w_3441_);
and (w_1347_, w_0841_, w_3104_);
or (w_2221_, w_2060_, w_1098_);
and (w_3516_, w_2615_, w_2325_);
or (w_1170_, w_2658_, w_0658_);
or (w_3058_, w_0390_, w_3216_);
and (out14[6], w_2087_, w_2347_);
or (w_0101_, w_2049_, w_2132_);
or (w_1761_, w_0878_, w_2856_);
or (w_3108_, w_3201_, w_0805_);
not (w_0371_, w_0090_);
and (w_2829_, w_2090_, w_0530_);
and (w_0210_, w_2509_, w_1905_);
or (w_2013_, w_1924_, w_1487_);
or (w_0035_, w_2206_, w_0416_);
or (w_3101_, w_1242_, w_1817_);
not (w_0422_, w_3451_);
or (w_2443_, in4[0], w_2994_);
and (w_0785_, w_1969_, w_0482_);
not (w_1536_, w_0161_);
or (w_1311_, w_0974_, w_2369_);
or (w_0076_, w_2581_, w_3364_);
or (w_2794_, out14[7], w_1849_);
not (w_2451_, in8[5]);
not (w_0640_, w_1267_);
not (w_1717_, w_2202_);
or (w_0961_, w_3199_, w_2114_);
or (w_0228_, w_0305_, w_1431_);
not (w_3142_, w_0624_);
and (w_3514_, w_2671_, w_3441_);
and (w_1326_, w_2197_, w_1064_);
and (out22[0], w_1036_, w_1180_);
and (w_0267_, w_1374_, w_0775_);
not (w_2037_, w_0829_);
not (w_1286_, in1[3]);
and (out6[5], w_3497_, w_0658_);
and (w_1595_, in3[4], w_2699_);
and (w_0913_, w_1429_, w_2073_);
not (w_0751_, w_0933_);
or (w_0408_, w_2559_, w_0630_);
and (w_0798_, in6[1], w_0872_);
not (w_0456_, w_3218_);
not (w_0554_, w_2248_);
or (w_0742_, w_2131_, w_2672_);
and (w_2572_, w_1466_, w_1030_);
or (w_1046_, w_3006_, w_0309_);
and (w_2632_, w_0387_, w_1873_);
and (w_0737_, w_3491_, w_0702_);
or (w_0349_, w_2435_, w_2519_);
not (w_2110_, w_3120_);
or (w_0292_, w_3253_, w_0518_);
and (w_3460_, w_2333_, w_2916_);
or (w_2285_, w_2788_, w_0142_);
or (w_0664_, w_0671_, w_2803_);
or (w_0181_, w_3408_, w_3169_);
or (w_3118_, w_2619_, w_2771_);
or (w_2589_, w_0601_, w_0710_);
or (w_1729_, out13[7], w_0929_);
or (w_0727_, w_2362_, w_1714_);
or (out23[1], w_2759_, w_0853_);
and (w_2515_, in7[5], w_1571_);
not (w_2087_, w_2660_);
or (w_2058_, in12[0], w_3160_);
not (w_2704_, w_2388_);
or (w_2297_, w_2370_, w_1307_);
and (w_1205_, w_2676_, w_3027_);
and (w_2712_, w_0149_, w_2148_);
and (w_1352_, w_1122_, w_1839_);
or (w_3469_, w_1719_, w_2580_);
and (w_0949_, w_2618_, w_0121_);
not (w_2400_, w_2906_);
not (w_3084_, w_2171_);
not (w_0736_, w_2100_);
and (out24[1], w_1630_, w_2133_);
or (w_2125_, w_1536_, w_1266_);
or (w_3143_, w_1141_, w_3183_);
not (w_3385_, w_0712_);
or (w_0060_, w_0824_, w_0950_);
and (w_0276_, w_1114_, w_1115_);
or (w_0838_, in12[1], w_0777_);
and (w_2028_, w_3218_, w_0658_);
or (w_2177_, w_3388_, w_0718_);
and (w_1240_, w_0749_, w_1567_);
or (w_3358_, w_3465_, w_2696_);
or (w_2928_, w_1108_, w_3319_);
and (w_2566_, w_0042_, w_2731_);
or (w_3092_, w_0265_, w_1951_);
and (w_1897_, w_0041_, w_2303_);
not (w_1258_, w_0859_);
or (w_2913_, w_3227_, w_2306_);
or (w_1525_, w_1666_, w_3050_);
or (w_3487_, w_1622_, w_2996_);
or (w_1565_, w_2393_, w_3042_);
or (w_1998_, w_1474_, w_1495_);
not (w_0032_, w_0137_);
not (w_0809_, in14[1]);
and (w_0609_, w_1535_, w_3222_);
and (w_2642_, w_0416_, w_3292_);
or (w_0723_, w_1535_, w_1737_);
or (w_1265_, in7[5], w_2800_);
and (w_0743_, in9[4], in10[0]);
and (w_0596_, w_2935_, w_1030_);
or (w_0475_, in5[0], w_2914_);
or (w_3113_, w_1359_, w_2798_);
and (w_3408_, in8[4], w_3184_);
or (w_0004_, w_0772_, w_1189_);
not (w_2941_, w_1304_);
or (w_0447_, w_3295_, w_0625_);
and (w_1047_, w_2184_, w_3380_);
or (w_0756_, w_2340_, w_3521_);
or (w_0778_, w_2009_, w_3269_);
and (w_0559_, w_1978_, w_2528_);
or (w_0190_, w_0913_, w_2472_);
and (w_0336_, w_1589_, w_2684_);
or (w_1051_, w_1719_, w_2959_);
or (w_1741_, in9[2], in10[2]);
or (w_2078_, w_1242_, w_2436_);
not (w_2290_, w_3393_);
and (w_0204_, w_0452_, w_1516_);
and (w_3449_, w_0909_, w_0098_);
or (w_2908_, w_0009_, w_2379_);
or (w_0011_, w_0143_, w_3071_);
and (w_2389_, w_3352_, w_3426_);
not (w_0387_, in7[1]);
and (w_1174_, w_0151_, w_2554_);
or (w_3154_, w_1420_, w_1489_);
or (w_3424_, w_3405_, w_2570_);
or (w_2693_, w_2516_, w_3102_);
and (w_1961_, in9[7], in10[7]);
and (w_2818_, w_2716_, w_1453_);
or (w_0775_, in9[6], in10[6]);
and (out13[2], w_2050_, w_3117_);
or (w_0947_, w_1246_, w_2068_);
and (w_3446_, w_0285_, w_0954_);
or (w_1268_, out13[7], w_0342_);
not (w_0039_, w_0084_);
or (w_0167_, w_2140_, w_2691_);
or (w_0314_, w_0258_, w_1988_);
and (w_0308_, w_2810_, out16[7]);
not (w_2621_, w_1009_);
or (w_3036_, w_1468_, w_0979_);
or (w_3312_, w_1041_, w_0134_);
and (w_0259_, w_0457_, w_1412_);
and (w_3525_, w_0045_, w_2296_);
or (w_0957_, in16[4], w_3132_);
and (w_2815_, w_2735_, w_2458_);
and (w_2924_, w_0669_, w_1535_);
not (w_1490_, w_1693_);
not (w_2713_, w_2858_);
or (w_1644_, w_1194_, w_0376_);
and (w_1510_, w_1045_, w_2407_);
or (w_0068_, in6[3], w_3483_);
not (w_3252_, w_2705_);
and (w_2960_, w_3501_, w_3287_);
or (w_3200_, w_0916_, w_1508_);
and (w_3078_, w_2963_, w_1164_);
and (w_3208_, in6[1], in5[0]);
and (w_2830_, w_0657_, w_1004_);
or (w_3102_, w_1417_, w_2029_);
and (w_2197_, w_1716_, w_2610_);
and (w_3401_, w_1227_, w_2208_);
and (w_1629_, w_0639_, w_0505_);
or (w_1895_, w_0987_, w_2113_);
not (w_2902_, w_0706_);
or (w_1538_, w_2207_, w_2674_);
or (w_0206_, w_1978_, w_2528_);
and (w_2355_, w_2429_, w_2018_);
and (w_2100_, w_1551_, w_3290_);
and (w_1851_, w_3237_, w_1518_);
not (w_1628_, in3[4]);
and (w_2961_, w_0141_, w_1517_);
not (w_3289_, w_0404_);
or (w_3406_, w_1670_, w_1493_);
or (w_2858_, w_3390_, w_3069_);
and (w_0283_, w_1320_, w_3337_);
and (w_0875_, w_2228_, w_0828_);
not (w_2426_, w_3361_);
or (w_0122_, w_1983_, w_1730_);
and (w_1154_, w_1871_, w_1018_);
and (w_1881_, w_3433_, w_2799_);
and (w_0517_, w_1459_, w_2084_);
or (out19[5], w_3470_, w_3110_);
and (w_1919_, w_0429_, w_0075_);
or (w_3112_, w_2077_, w_1350_);
or (w_3488_, w_3194_, w_2871_);
or (w_2213_, w_3302_, w_1335_);
or (w_3136_, w_1983_, w_0426_);
and (w_2951_, w_0322_, w_2517_);
or (w_1646_, in8[5], w_1076_);
and (w_0125_, w_2990_, w_1029_);
or (w_1549_, w_2476_, w_2142_);
or (w_1740_, w_2873_, w_2439_);
or (w_1139_, w_3331_, w_0822_);
or (w_1985_, w_2281_, w_0433_);
or (w_0698_, w_2000_, w_0118_);
not (w_1204_, w_3082_);
or (w_3273_, w_3156_, w_2628_);
not (w_1848_, w_2204_);
and (w_1997_, w_2086_, w_2371_);
or (w_1816_, w_3091_, w_2971_);
or (w_3321_, in15[1], w_1213_);
not (w_1489_, w_2994_);
and (out22[5], w_1438_, w_1749_);
not (w_0264_, w_3453_);
and (w_0436_, w_2942_, w_2781_);
or (w_3213_, w_0456_, w_3088_);
or (w_2616_, w_2226_, w_1179_);
or (w_3477_, w_3519_, w_3478_);
or (w_1307_, w_2479_, w_2205_);
not (w_1082_, w_3208_);
and (w_0010_, in5[0], w_2914_);
or (w_1363_, w_0748_, w_3496_);
not (w_0459_, w_1382_);
and (w_2029_, w_3095_, w_2657_);
not (w_2366_, in15[1]);
not (w_3248_, w_0217_);
or (w_0454_, w_0963_, w_1424_);
not (w_0865_, in14[4]);
not (w_1006_, w_1880_);
and (w_0695_, w_1673_, w_0712_);
and (w_2545_, w_1910_, w_1103_);
and (w_1065_, w_2409_, w_1458_);
or (w_0962_, w_3405_, w_0601_);
or (w_3524_, w_3218_, w_0658_);
or (w_0261_, w_1320_, w_0659_);
not (w_1269_, w_1635_);
not (w_0221_, w_1842_);
and (w_3122_, w_0888_, w_2293_);
and (w_3508_, w_2416_, w_2625_);
and (w_0566_, w_1655_, w_0171_);
and (w_1930_, w_0641_, w_2475_);
and (w_0374_, w_3492_, w_0512_);
and (w_3259_, w_2589_, w_1564_);
or (w_2341_, w_3493_, w_2026_);
or (w_1189_, w_0875_, w_2001_);
or (w_2991_, w_3141_, w_0502_);
not (w_1768_, w_0871_);
or (w_0280_, w_1714_, w_0747_);
or (w_2165_, w_0322_, w_2153_);
not (w_0665_, w_2304_);
or (w_0069_, w_0790_, w_0599_);
not (w_1906_, w_1836_);
or (w_3074_, w_0809_, w_2912_);
and (w_1447_, w_0365_, w_1886_);
and (w_1295_, w_0942_, w_0060_);
and (w_2264_, w_2042_, w_2276_);
or (w_1049_, w_2954_, w_1980_);
not (w_3222_, w_3292_);
or (w_1769_, w_2544_, w_1755_);
or (w_2303_, w_1570_, w_3457_);
or (w_2372_, w_0402_, w_2294_);
or (w_1931_, w_3268_, w_1327_);
not (w_3164_, w_3157_);
or (w_0658_, w_0057_, w_1283_);
or (w_2727_, in6[4], in5[3]);
or (w_2071_, w_3186_, w_0647_);
or (w_2997_, w_2566_, w_0046_);
or (w_2876_, w_1173_, w_1779_);
or (w_2765_, w_3264_, w_2301_);
or (w_1614_, w_2883_, w_1754_);
not (w_2049_, out13[7]);
or (w_3021_, w_1203_, w_3411_);
and (w_0250_, w_0312_, w_2399_);
or (w_1977_, w_3146_, w_1650_);
and (w_2496_, in1[0], in2[1]);
and (w_0831_, in11[6], w_1465_);
or (w_2311_, w_3308_, w_0054_);
or (w_0923_, w_1290_, w_0769_);
not (w_2159_, w_0259_);
and (w_0419_, w_2440_, w_2693_);
or (w_0510_, in12[5], w_0740_);
not (w_0432_, w_2279_);
or (w_3430_, w_1758_, w_2902_);
not (w_3319_, w_2041_);
and (w_3519_, w_3412_, w_0804_);
or (w_1624_, w_0019_, w_1836_);
or (w_1532_, w_0649_, w_0470_);
or (w_0290_, w_1648_, w_0918_);
and (w_2047_, w_2738_, w_1721_);
or (w_2720_, w_1209_, w_1705_);
and (w_1453_, w_2760_, w_2834_);
or (w_1023_, w_1326_, w_3414_);
not (w_0545_, w_3503_);
and (w_2591_, w_2773_, w_1050_);
and (w_2842_, w_3403_, w_0206_);
or (w_0830_, w_0006_, w_3513_);
not (w_1876_, w_1949_);
not (w_0256_, w_0716_);
or (w_1341_, w_0044_, w_1454_);
not (w_1853_, w_2064_);
not (w_2931_, w_0839_);
or (w_1822_, w_3209_, w_1686_);
and (w_3232_, w_1553_, w_0043_);
or (w_0682_, w_1183_, w_2783_);
or (w_2042_, w_1275_, w_3292_);
not (w_3338_, w_0984_);
or (w_2195_, w_0783_, w_0574_);
or (w_2217_, w_1141_, w_3492_);
or (w_1803_, w_2051_, w_1565_);
and (w_2660_, w_3058_, w_1148_);
and (w_0783_, w_2339_, w_3018_);
or (w_2527_, w_1691_, w_2709_);
or (w_0709_, w_2677_, w_3221_);
or (w_2937_, w_0032_, w_2286_);
and (w_1574_, w_3157_, w_2287_);
and (w_1755_, w_0329_, w_0642_);
or (w_1200_, w_1246_, w_2141_);
not (w_0464_, w_1811_);
and (w_2233_, in5[5], w_0975_);
or (w_3383_, w_1156_, w_3272_);
not (w_1374_, w_2364_);
or (w_2888_, w_1111_, w_1798_);
or (w_1135_, w_1000_, w_0663_);
not (w_3440_, out16[2]);
or (w_2231_, w_3328_, w_3183_);
and (w_0509_, w_3527_, w_0951_);
and (w_1213_, w_1394_, w_0882_);
not (w_0987_, w_1690_);
and (w_2331_, w_0074_, w_2403_);
not (w_1712_, w_0078_);
or (w_1445_, w_3487_, w_1126_);
or (w_3063_, w_2933_, w_1950_);
and (w_2918_, in4[2], w_2863_);
or (w_1656_, w_2593_, w_1790_);
not (w_0741_, w_3244_);
and (w_2907_, w_3506_, w_1584_);
or (w_1767_, w_1586_, w_2290_);
and (w_0095_, w_2213_, w_2973_);
and (w_3493_, w_2353_, w_0065_);
and (w_0750_, w_1719_, w_0421_);
and (out1[4], w_1051_, w_2681_);
or (out15[7], w_1953_, w_3281_);
or (w_1613_, w_3192_, w_1201_);
and (w_1659_, w_0130_, w_2002_);
or (w_0452_, w_0339_, w_0948_);
not (w_1569_, w_2800_);
and (w_0208_, w_0511_, w_1470_);
not (w_3111_, w_3191_);
or (w_1687_, w_1823_, w_1254_);
and (w_2751_, w_1640_, w_2886_);
or (w_2444_, w_2091_, w_2932_);
and (w_0080_, w_3426_, w_2901_);
not (w_1995_, w_1295_);
and (w_1310_, w_2944_, w_3389_);
and (w_2903_, w_0790_, w_3501_);
and (w_0732_, w_2194_, w_2438_);
not (w_1331_, w_0592_);
or (w_0749_, w_1501_, w_1706_);
or (w_0992_, w_2576_, w_2720_);
not (w_1630_, w_1100_);
or (w_2461_, w_0001_, w_3376_);
or (w_0149_, w_3293_, w_2510_);
not (w_0383_, w_3229_);
not (w_2336_, w_1861_);
not (w_1008_, w_0919_);
not (w_1570_, w_0725_);
or (w_2420_, w_1644_, w_3528_);
not (w_2276_, w_0473_);
and (w_1040_, w_1224_, w_2529_);
and (w_2569_, w_1176_, w_0179_);
not (w_1929_, w_2179_);
or (w_3018_, w_1746_, w_0753_);
not (w_0340_, in1[1]);
or (w_1294_, w_1541_, w_3162_);
and (w_3331_, in3[3], w_2892_);
not (w_0199_, w_3428_);
and (w_1002_, w_3368_, w_2224_);
and (w_1917_, w_2736_, w_3440_);
or (w_1171_, w_0618_, w_2502_);
or (w_2964_, w_0237_, w_2139_);
or (w_0860_, w_0579_, w_2604_);
or (w_2486_, in6[4], w_0526_);
or (w_1976_, w_0271_, w_3297_);
and (w_2437_, w_3417_, w_2861_);
or (w_1208_, w_0501_, w_2387_);
not (w_2917_, w_0619_);
not (w_0514_, in13[1]);
and (w_1763_, in9[2], in10[2]);
and (w_2008_, w_2131_, w_3060_);
or (w_2395_, w_1084_, w_0776_);
or (w_3100_, w_2873_, w_0717_);
and (w_0416_, w_1569_, w_2906_);
not (w_1469_, w_3509_);
or (w_3056_, w_0862_, w_1396_);
or (w_0702_, w_2718_, w_0675_);
and (w_2005_, w_0696_, w_0953_);
and (w_0347_, w_1535_, w_1737_);
and (w_2163_, w_2214_, w_2929_);
or (w_3288_, w_0852_, w_2003_);
or (out19[0], w_0601_, w_3394_);
or (w_1444_, w_2339_, w_3018_);
and (w_0470_, w_1771_, w_0799_);
or (w_1677_, w_0804_, w_0658_);
or (w_0650_, w_3333_, w_3195_);
and (w_2708_, w_1676_, w_2288_);
or (w_3235_, w_0804_, w_3426_);
not (w_3203_, in5[4]);
and (w_1751_, w_0458_, w_2829_);
or (w_2756_, w_0125_, w_3046_);
and (w_2665_, in15[2], w_2176_);
and (w_3028_, w_2444_, w_3235_);
or (w_1131_, w_3189_, w_1979_);
and (w_0505_, w_0988_, w_0093_);
or (w_2672_, w_1848_, w_2768_);
not (w_1649_, w_3457_);
or (w_1001_, w_2717_, w_3059_);
not (w_0325_, w_0193_);
not (w_3009_, w_1832_);
or (w_2488_, w_1474_, w_3060_);
and (w_0014_, w_0472_, w_2821_);
or (w_0391_, in12[1], w_2943_);
or (w_0360_, w_2511_, w_3399_);
and (w_0621_, w_2172_, w_2897_);
and (w_1620_, w_1393_, w_2614_);
and (out10[0], w_0079_, w_3317_);
or (w_1904_, w_1521_, w_2653_);
not (w_2667_, w_2153_);
or (w_1407_, w_2578_, w_0604_);
or (w_2570_, w_0265_, w_0459_);
and (w_3053_, w_2196_, w_0400_);
or (w_0321_, w_1547_, w_1587_);
and (w_2344_, w_1429_, w_1535_);
or (w_1794_, w_2646_, w_1199_);
and (w_0768_, in7[5], w_2800_);
and (w_3310_, w_2027_, w_1153_);
or (w_0836_, w_1436_, w_1531_);
and (w_3156_, w_3297_, w_0760_);
endmodule

module sub_module3(
    input wire [1:0] in1,
    input wire [1:0] in2,
    input wire [1:0] in3,
    input wire [1:0] in4,
    input wire [1:0] in5,
    input wire [1:0] in6,
    input wire [1:0] in7,
    input wire [1:0] in8,
    input wire [1:0] in9,
    input wire [1:0] in10,
    input wire [1:0] in11,
    input wire [1:0] in12,
    input wire [1:0] in13,
    input wire [1:0] in14,
    input wire [1:0] in15,
    output wire out1,
    output wire out2,
    output wire out3,
    output wire out4,
    output wire out5,
    output wire out6,
    output wire out7,
    output wire out8,
    output wire out9,
    output wire out10,
    output wire out11,
    output wire out12,
    output wire out13,
    output wire out14,
    output wire out15
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
or (w_0238_, w_0117_, w_0708_);
or (w_0129_, w_0581_, w_0118_);
or (w_0488_, w_0212_, w_0136_);
and (w_0019_, w_0510_, w_0344_);
or (w_0174_, w_0243_, w_0025_);
and (w_0137_, w_0293_, w_0421_);
and (w_0136_, w_0106_, w_0363_);
and (w_0446_, w_0133_, w_0447_);
and (w_0278_, w_0581_, w_0173_);
or (w_0101_, in15[0], w_0475_);
or (w_0031_, w_0720_, w_0185_);
and (w_0110_, w_0545_, w_0513_);
or (w_0038_, w_0406_, w_0206_);
or (out13, w_0536_, w_0357_);
and (w_0145_, w_0836_, w_0115_);
and (w_0536_, in15[1], w_0242_);
not (w_0248_, in9[0]);
or (w_0834_, w_0191_, w_0201_);
and (w_0618_, in13[0], in14[0]);
or (w_0065_, w_0655_, w_0779_);
or (w_0023_, in3[1], in4[1]);
or (w_0253_, w_0103_, w_0511_);
or (w_0099_, w_0631_, w_0815_);
or (w_0763_, w_0764_, w_0317_);
and (w_0349_, w_0599_, w_0839_);
and (w_0230_, w_0098_, w_0020_);
and (w_0184_, w_0051_, w_0574_);
and (w_0704_, w_0284_, w_0630_);
and (w_0530_, w_0675_, w_0105_);
and (w_0608_, in15[0], w_0475_);
or (w_0437_, w_0726_, w_0257_);
or (w_0805_, w_0311_, w_0075_);
or (w_0379_, w_0205_, w_0692_);
and (w_0443_, w_0413_, w_0681_);
and (w_0382_, w_0755_, w_0609_);
and (w_0594_, w_0282_, w_0687_);
and (w_0378_, w_0599_, w_0156_);
and (w_0517_, w_0098_, w_0165_);
and (w_0575_, w_0581_, w_0523_);
not (w_0183_, w_0369_);
or (w_0831_, w_0375_, w_0312_);
or (w_0263_, w_0388_, w_0481_);
or (w_0296_, w_0450_, w_0265_);
or (w_0641_, w_0396_, w_0629_);
and (w_0114_, w_0004_, w_0785_);
and (w_0152_, in15[1], w_0181_);
or (w_0005_, w_0598_, w_0363_);
and (w_0794_, w_0237_, w_0486_);
or (w_0791_, in7[0], in8[0]);
or (w_0541_, w_0110_, w_0594_);
or (w_0167_, w_0210_, w_0488_);
and (w_0445_, w_0507_, w_0689_);
or (w_0532_, in15[0], w_0547_);
and (w_0607_, w_0816_, w_0010_);
and (w_0728_, w_0063_, w_0766_);
or (out5, w_0427_, w_0462_);
and (w_0163_, w_0734_, w_0826_);
and (w_0160_, w_0236_, w_0390_);
or (w_0073_, w_0081_, w_0186_);
not (w_0341_, in9[1]);
or (w_0664_, w_0374_, w_0058_);
and (w_0388_, w_0432_, w_0549_);
and (w_0175_, w_0091_, w_0062_);
or (w_0843_, w_0033_, w_0081_);
or (w_0472_, w_0180_, w_0634_);
or (w_0074_, w_0651_, w_0016_);
and (w_0474_, w_0233_, w_0698_);
and (w_0100_, w_0192_, w_0470_);
not (w_0318_, w_0486_);
and (w_0552_, w_0081_, w_0186_);
and (w_0537_, w_0307_, w_0483_);
or (w_0280_, w_0618_, w_0755_);
or (w_0747_, w_0461_, w_0684_);
or (w_0813_, w_0652_, w_0485_);
and (w_0053_, in5[0], in6[1]);
or (w_0688_, w_0425_, w_0490_);
or (w_0182_, w_0411_, w_0750_);
or (w_0094_, w_0125_, w_0497_);
and (w_0035_, w_0153_, w_0645_);
and (w_0390_, w_0662_, w_0006_);
or (w_0311_, w_0772_, w_0083_);
or (w_0106_, in1[1], in2[0]);
and (w_0660_, w_0583_, w_0041_);
and (w_0372_, w_0093_, w_0633_);
or (w_0554_, w_0027_, w_0585_);
or (w_0557_, w_0192_, w_0801_);
and (w_0146_, w_0581_, w_0632_);
and (w_0565_, w_0791_, w_0225_);
or (w_0696_, w_0776_, w_0321_);
and (w_0701_, w_0730_, w_0731_);
or (w_0307_, w_0336_, w_0229_);
and (w_0543_, w_0034_, w_0420_);
and (w_0356_, w_0473_, w_0051_);
and (w_0141_, w_0149_, w_0397_);
or (w_0143_, w_0572_, w_0019_);
and (w_0376_, w_0417_, w_0559_);
and (w_0239_, w_0728_, w_0778_);
and (w_0133_, w_0341_, w_0218_);
or (w_0746_, w_0002_, w_0042_);
not (w_0322_, w_0005_);
and (w_0267_, w_0098_, w_0148_);
or (w_0473_, w_0219_, w_0268_);
or (out11, w_0347_, w_0517_);
and (w_0485_, w_0237_, w_0624_);
and (w_0774_, w_0733_, w_0721_);
and (w_0459_, w_0634_, w_0485_);
and (w_0273_, w_0568_, w_0659_);
or (w_0513_, w_0079_, w_0365_);
or (w_0758_, in15[0], w_0767_);
or (w_0172_, w_0329_, w_0601_);
or (w_0144_, w_0034_, w_0420_);
and (w_0034_, w_0773_, w_0843_);
or (w_0015_, w_0040_, w_0018_);
and (w_0040_, w_0304_, w_0476_);
not (w_0218_, in10[0]);
and (w_0203_, w_0426_, w_0564_);
and (w_0544_, w_0129_, w_0335_);
and (w_0112_, w_0779_, w_0705_);
and (w_0438_, w_0255_, w_0338_);
or (w_0394_, w_0842_, w_0759_);
and (w_0374_, in15[0], w_0137_);
or (w_0115_, w_0383_, w_0071_);
not (w_0084_, w_0457_);
or (w_0085_, w_0113_, w_0403_);
or (w_0449_, w_0409_, w_0479_);
and (w_0285_, w_0098_, w_0695_);
and (w_0694_, w_0052_, w_0360_);
and (w_0605_, w_0830_, w_0508_);
or (w_0600_, w_0605_, w_0149_);
or (w_0018_, w_0649_, w_0184_);
not (w_0776_, in7[0]);
and (w_0180_, in2[1], in1[0]);
or (w_0503_, w_0613_, w_0059_);
and (w_0012_, w_0286_, w_0686_);
or (w_0419_, w_0003_, w_0453_);
or (w_0785_, w_0237_, w_0486_);
and (w_0482_, in15[1], w_0544_);
or (w_0646_, w_0478_, w_0080_);
or (w_0313_, w_0736_, w_0359_);
or (w_0000_, w_0032_, w_0777_);
and (w_0679_, w_0605_, w_0149_);
and (w_0745_, w_0658_, w_0541_);
and (w_0255_, w_0800_, w_0245_);
or (out8, w_0152_, w_0230_);
and (w_0279_, w_0065_, w_0249_);
and (w_0418_, in15[1], w_0484_);
and (w_0214_, w_0686_, w_0619_);
or (w_0705_, in9[0], in10[0]);
or (w_0609_, w_0710_, w_0195_);
and (w_0147_, w_0210_, w_0488_);
and (w_0559_, w_0558_, w_0094_);
and (w_0397_, w_0188_, w_0835_);
and (w_0616_, in15[0], w_0767_);
and (w_0201_, w_0401_, w_0323_);
or (w_0309_, w_0307_, w_0483_);
or (w_0346_, w_0781_, w_0472_);
and (w_0261_, w_0092_, w_0566_);
or (w_0006_, w_0310_, w_0833_);
or (w_0158_, w_0550_, w_0610_);
or (w_0844_, w_0368_, w_0788_);
or (w_0348_, w_0837_, w_0337_);
or (w_0533_, w_0214_, w_0459_);
or (w_0275_, w_0069_, w_0408_);
or (w_0663_, w_0023_, w_0652_);
and (w_0639_, w_0598_, w_0425_);
or (w_0092_, w_0581_, w_0489_);
or (w_0235_, w_0097_, w_0100_);
and (w_0332_, in15[0], w_0824_);
and (w_0837_, w_0279_, w_0496_);
or (w_0693_, w_0570_, w_0379_);
and (w_0398_, w_0023_, w_0652_);
or (w_0060_, in15[0], w_0491_);
or (w_0272_, w_0755_, w_0609_);
and (w_0260_, w_0703_, w_0618_);
or (w_0042_, w_0552_, w_0745_);
and (w_0752_, w_0673_, w_0172_);
or (w_0191_, in13[0], in14[0]);
and (w_0534_, w_0568_, w_0298_);
and (w_0281_, in1[1], in2[0]);
and (w_0789_, w_0098_, w_0209_);
not (w_0321_, in8[1]);
or (w_0784_, w_0621_, w_0057_);
and (w_0016_, w_0263_, w_0002_);
and (w_0242_, w_0270_, w_0101_);
and (w_0571_, w_0422_, w_0248_);
and (w_0519_, w_0460_, w_0740_);
and (w_0560_, w_0098_, w_0664_);
or (w_0464_, w_0460_, w_0287_);
or (w_0192_, w_0088_, w_0766_);
and (w_0125_, w_0841_, w_0393_);
and (w_0294_, w_0807_, w_0300_);
or (w_0416_, w_0282_, w_0687_);
or (w_0807_, w_0836_, w_0115_);
and (w_0177_, w_0168_, w_0791_);
or (w_0623_, w_0164_, w_0011_);
not (w_0258_, in4[1]);
or (w_0779_, w_0248_, w_0218_);
and (w_0547_, w_0648_, w_0194_);
or (w_0236_, in11[0], in12[1]);
and (w_0743_, w_0032_, w_0777_);
and (w_0371_, w_0167_, w_0592_);
or (w_0373_, w_0236_, w_0339_);
and (w_0441_, w_0563_, w_0056_);
and (w_0027_, w_0341_, w_0422_);
and (w_0637_, w_0577_, w_0676_);
and (w_0276_, w_0098_, w_0277_);
or (w_0165_, w_0244_, w_0223_);
and (w_0402_, in15[0], w_0683_);
and (w_0155_, w_0440_, w_0790_);
not (w_0107_, w_0705_);
and (w_0302_, w_0206_, w_0619_);
and (w_0257_, w_0425_, w_0444_);
or (w_0298_, w_0505_, w_0786_);
or (w_0835_, w_0791_, w_0225_);
or (w_0249_, w_0660_, w_0003_);
and (w_0468_, w_0423_, w_0448_);
and (w_0139_, w_0015_, w_0246_);
or (w_0838_, w_0128_, w_0449_);
and (w_0440_, in14[0], in13[1]);
and (w_0720_, in12[0], in11[1]);
and (w_0122_, w_0385_, w_0626_);
and (w_0606_, w_0174_, w_0182_);
and (w_0083_, w_0021_, w_0658_);
or (w_0454_, w_0106_, w_0363_);
or (w_0264_, w_0599_, w_0839_);
and (w_0516_, w_0125_, w_0320_);
or (w_0709_, in10[1], in9[0]);
and (w_0069_, w_0492_, w_0757_);
and (w_0024_, w_0098_, w_0756_);
and (w_0615_, w_0831_, w_0133_);
or (w_0131_, w_0204_, w_0108_);
and (w_0665_, w_0327_, w_0734_);
or (w_0659_, w_0160_, w_0438_);
and (w_0025_, w_0582_, w_0650_);
and (w_0749_, w_0581_, w_0118_);
or (w_0632_, w_0260_, w_0606_);
or (w_0514_, in15[0], w_0207_);
and (w_0748_, w_0673_, w_0158_);
or (w_0523_, w_0519_, w_0273_);
not (w_0304_, in12[0]);
and (w_0790_, w_0802_, w_0130_);
or (w_0148_, w_0332_, w_0077_);
and (w_0611_, in9[1], in10[1]);
or (w_0699_, w_0410_, w_0540_);
or (w_0727_, w_0274_, w_0804_);
not (w_0810_, w_0154_);
and (w_0685_, w_0038_, w_0663_);
or (w_0447_, w_0565_, w_0553_);
and (w_0226_, w_0103_, w_0511_);
and (w_0392_, w_0655_, w_0779_);
and (w_0667_, in15[1], w_0261_);
or (w_0228_, w_0324_, w_0269_);
or (w_0598_, in1[1], in2[1]);
or (w_0051_, w_0027_, w_0611_);
or (w_0224_, w_0616_, w_0043_);
or (w_0385_, w_0728_, w_0533_);
or (w_0179_, w_0068_, w_0429_);
and (w_0569_, w_0164_, w_0011_);
and (w_0803_, w_0836_, w_0149_);
or (w_0756_, w_0289_, w_0501_);
and (w_0478_, w_0827_, w_0321_);
and (w_0377_, w_0281_, w_0358_);
and (w_0452_, w_0000_, w_0031_);
and (w_0409_, w_0842_, w_0759_);
and (w_0432_, w_0044_, w_0189_);
or (w_0190_, w_0568_, w_0659_);
and (w_0715_, w_0776_, w_0321_);
or (w_0011_, w_0794_, w_0713_);
or (w_0592_, w_0455_, w_0315_);
or (w_0271_, in7[0], in8[1]);
and (w_0268_, w_0844_, w_0510_);
or (w_0799_, w_0351_, w_0234_);
and (w_0355_, in15[0], w_0424_);
and (w_0584_, w_0652_, w_0485_);
and (w_0043_, w_0581_, w_0763_);
or (w_0002_, w_0075_, w_0440_);
and (w_0353_, in10[1], in9[0]);
and (w_0059_, w_0128_, w_0449_);
and (w_0369_, in7[0], in8[0]);
or (w_0384_, w_0504_, w_0506_);
not (w_0098_, in15[1]);
and (w_0484_, w_0671_, w_0532_);
and (w_0590_, w_0135_, w_0697_);
and (w_0220_, in15[1], w_0530_);
not (w_0713_, w_0785_);
or (w_0451_, w_0562_, w_0162_);
and (w_0771_, w_0714_, w_0758_);
or (w_0426_, w_0614_, w_0334_);
or (w_0757_, w_0556_, w_0048_);
and (w_0540_, w_0493_, w_0045_);
or (w_0840_, w_0334_, w_0222_);
or (w_0714_, w_0581_, w_0763_);
and (w_0457_, w_0197_, w_0106_);
or (w_0690_, w_0543_, w_0333_);
and (w_0809_, in6[0], in5[1]);
and (w_0760_, w_0587_, w_0466_);
or (w_0362_, w_0473_, w_0051_);
or (w_0173_, w_0017_, w_0217_);
and (w_0580_, w_0787_, w_0088_);
and (w_0326_, w_0812_, w_0478_);
or (w_0502_, w_0581_, w_0124_);
and (w_0297_, in15[0], w_0480_);
and (w_0181_, w_0216_, w_0292_);
and (w_0256_, w_0455_, w_0315_);
or (w_0266_, w_0665_, w_0326_);
or (w_0630_, w_0492_, w_0757_);
and (w_0219_, w_0647_, w_0504_);
or (w_0579_, w_0299_, w_0035_);
or (w_0833_, w_0256_, w_0147_);
and (w_0357_, w_0098_, w_0029_);
and (w_0460_, in14[1], in13[1]);
not (w_0653_, in3[1]);
and (w_0327_, w_0309_, w_0251_);
and (w_0628_, in15[1], w_0372_);
or (w_0001_, w_0468_, w_0829_);
and (w_0128_, w_0411_, w_0622_);
or (w_0563_, w_0153_, w_0306_);
and (w_0414_, w_0660_, w_0003_);
and (w_0247_, w_0098_, w_0717_);
and (w_0804_, w_0030_, w_0170_);
and (w_0677_, w_0391_, w_0701_);
and (w_0741_, w_0027_, w_0585_);
or (w_0246_, w_0161_, w_0591_);
not (w_0229_, w_0393_);
and (w_0310_, w_0709_, w_0718_);
or (w_0836_, w_0341_, w_0218_);
and (w_0829_, w_0121_, w_0211_);
or (w_0196_, w_0236_, w_0390_);
and (w_0825_, w_0036_, w_0729_);
or (w_0830_, w_0132_, w_0822_);
not (w_0680_, w_0657_);
and (w_0367_, w_0081_, w_0150_);
not (w_0622_, in14[1]);
and (w_0185_, w_0576_, w_0600_);
or (w_0662_, w_0798_, w_0371_);
or (w_0508_, w_0538_, w_0350_);
and (w_0078_, in15[1], w_0431_);
and (w_0111_, w_0562_, w_0162_);
or (w_0213_, w_0206_, w_0619_);
and (w_0627_, w_0032_, w_0161_);
and (w_0480_, w_0190_, w_0364_);
and (w_0733_, w_0204_, w_0192_);
not (w_0412_, w_0237_);
and (w_0316_, w_0728_, w_0301_);
or (w_0739_, w_0314_, w_0781_);
and (w_0490_, in1[0], in2[0]);
and (w_0113_, w_0589_, w_0275_);
or (w_0386_, w_0053_, w_0784_);
or (w_0157_, w_0571_, w_0579_);
and (w_0625_, w_0620_, w_0578_);
and (w_0716_, in15[1], w_0821_);
not (w_0004_, w_0794_);
or (w_0689_, w_0432_, w_0549_);
and (w_0080_, in7[1], in8[1]);
and (w_0221_, w_0098_, w_0224_);
or (w_0466_, w_0082_, w_0193_);
and (w_0193_, w_0425_, w_0012_);
not (w_0057_, w_0290_);
or (w_0797_, w_0589_, w_0128_);
or (w_0202_, w_0581_, w_0723_);
or (w_0216_, w_0581_, w_0173_);
or (w_0681_, w_0327_, w_0734_);
not (w_0088_, in5[1]);
and (w_0380_, in4[1], in3[0]);
and (w_0636_, w_0182_, w_0191_);
and (w_0475_, w_0272_, w_0834_);
or (w_0134_, w_0661_, w_0464_);
or (w_0130_, w_0081_, w_0150_);
or (w_0802_, w_0658_, w_0761_);
and (w_0842_, w_0782_, w_0419_);
and (w_0403_, w_0252_, w_0704_);
and (w_0821_, w_0711_, w_0387_);
or (w_0806_, w_0348_, w_0797_);
and (w_0231_, w_0625_, w_0702_);
and (w_0315_, w_0454_, w_0435_);
or (w_0200_, w_0297_, w_0575_);
or (w_0678_, w_0797_, w_0116_);
or (w_0455_, w_0226_, w_0070_);
or (w_0187_, w_0391_, w_0617_);
and (w_0410_, w_0068_, w_0429_);
and (w_0095_, w_0104_, w_0538_);
and (w_0642_, w_0098_, w_0238_);
or (w_0599_, w_0587_, w_0103_);
and (w_0710_, w_0759_, w_0294_);
or (w_0498_, w_0571_, w_0535_);
not (w_0211_, w_0611_);
or (w_0067_, w_0709_, w_0744_);
or (w_0370_, w_0841_, w_0670_);
and (w_0320_, w_0739_, w_0522_);
or (w_0072_, w_0391_, w_0028_);
or (w_0062_, in15[0], w_0050_);
or (w_0442_, w_0719_, w_0811_);
and (w_0365_, w_0271_, w_0803_);
and (w_0337_, w_0614_, w_0334_);
and (w_0090_, w_0581_, w_0085_);
or (w_0404_, w_0734_, w_0826_);
and (w_0644_, w_0391_, w_0028_);
and (w_0003_, in9[0], in10[0]);
or (w_0691_, w_0596_, w_0139_);
and (w_0755_, w_0411_, w_0750_);
or (w_0671_, w_0581_, w_0074_);
and (w_0826_, w_0526_, w_0140_);
and (w_0527_, w_0502_, w_0389_);
and (w_0786_, w_0334_, w_0222_);
or (w_0252_, w_0411_, w_0622_);
or (w_0056_, w_0080_, w_0122_);
and (w_0176_, w_0391_, w_0617_);
and (w_0077_, w_0581_, w_0489_);
or (out12, w_0340_, w_0022_);
and (w_0234_, w_0776_, w_0823_);
or (w_0524_, w_0715_, w_0436_);
and (w_0243_, w_0699_, w_0076_);
or (w_0511_, w_0234_, w_0369_);
or (w_0222_, w_0366_, w_0231_);
and (w_0070_, w_0192_, w_0801_);
and (w_0299_, w_0080_, w_0515_);
or (w_0640_, w_0603_, w_0208_);
or (out2, w_0716_, w_0247_);
or (w_0487_, w_0781_, w_0288_);
or (w_0086_, w_0322_, w_0198_);
or (w_0197_, in3[1], in4[0]);
not (w_0422_, in10[1]);
and (w_0726_, w_0781_, w_0288_);
or (w_0421_, w_0460_, w_0283_);
and (w_0406_, w_0653_, w_0258_);
and (w_0629_, w_0266_, w_0798_);
and (w_0469_, in15[0], w_0590_);
or (w_0269_, in6[0], in5[1]);
or (w_0525_, w_0625_, w_0702_);
or (w_0430_, w_0493_, w_0045_);
and (w_0028_, w_0813_, w_0213_);
and (w_0654_, w_0203_, w_0596_);
and (w_0055_, w_0169_, w_0754_);
and (w_0207_, w_0134_, w_0343_);
or (w_0673_, w_0580_, w_0809_);
or (w_0562_, w_0750_, w_0551_);
or (w_0127_, w_0733_, w_0685_);
or (w_0358_, w_0154_, w_0406_);
and (w_0643_, w_0709_, w_0744_);
and (w_0082_, w_0781_, w_0472_);
and (w_0303_, w_0486_, w_0154_);
and (w_0009_, w_0098_, w_0200_);
or (w_0135_, w_0252_, w_0704_);
and (w_0703_, w_0668_, w_0531_);
not (w_0166_, in4[0]);
not (w_0815_, in2[0]);
and (w_0081_, w_0171_, w_0700_);
and (w_0602_, w_0798_, w_0371_);
not (w_0551_, in13[1]);
or (w_0391_, in5[0], in6[1]);
or (w_0578_, w_0103_, w_0646_);
and (w_0491_, w_0548_, w_0573_);
and (w_0792_, w_0841_, w_0670_);
and (w_0651_, w_0445_, w_0407_);
or (out15, w_0259_, w_0221_);
and (w_0539_, w_0525_, w_0342_);
or (w_0751_, w_0781_, w_0099_);
or (w_0364_, w_0460_, w_0740_);
or (w_0153_, w_0827_, w_0321_);
not (w_0411_, in13[0]);
and (w_0395_, w_0039_, w_0060_);
or (w_0686_, in2[1], in1[0]);
or (out14, w_0220_, w_0009_);
and (w_0142_, w_0053_, w_0784_);
or (w_0583_, w_0819_, w_0132_);
and (w_0684_, w_0464_, w_0007_);
not (w_0500_, w_0722_);
or (w_0338_, w_0762_, w_0602_);
or (w_0542_, w_0055_, w_0607_);
and (w_0649_, w_0829_, w_0325_);
and (w_0538_, w_0271_, w_0696_);
or (w_0041_, w_0104_, w_0538_);
and (w_0505_, w_0496_, w_0539_);
or (w_0564_, w_0279_, w_0496_);
and (w_0458_, w_0661_, w_0464_);
or (w_0387_, in15[0], w_0381_);
not (w_0400_, w_0621_);
and (w_0259_, in15[1], w_0771_);
or (w_0399_, w_0599_, w_0156_);
or (w_0351_, w_0774_, w_0349_);
or (w_0595_, w_0496_, w_0539_);
or (w_0161_, in12[0], in11[1]);
and (w_0408_, w_0330_, w_0291_);
or (w_0029_, w_0608_, w_0199_);
and (w_0610_, w_0428_, w_0444_);
and (w_0839_, w_0722_, w_0037_);
and (w_0549_, in11[0], in12[1]);
and (w_0014_, w_0658_, w_0761_);
and (w_0736_, w_0003_, w_0453_);
and (w_0045_, w_0187_, w_0178_);
or (w_0510_, w_0823_, w_0827_);
or (w_0778_, w_0302_, w_0584_);
and (w_0650_, w_0067_, w_0498_);
and (w_0381_, w_0805_, w_0144_);
and (w_0151_, w_0456_, w_0073_);
or (w_0323_, w_0759_, w_0294_);
or (w_0735_, w_0215_, w_0832_);
or (w_0576_, w_0831_, w_0133_);
and (w_0075_, w_0750_, w_0551_);
or (w_0044_, w_0266_, w_0798_);
and (w_0103_, in5[1], in6[1]);
or (w_0162_, w_0367_, w_0014_);
and (w_0596_, w_0252_, w_0603_);
or (w_0188_, w_0234_, w_0593_);
and (w_0529_, w_0810_, w_0023_);
or (w_0574_, w_0163_, w_0467_);
and (w_0767_, w_0678_, w_0691_);
and (w_0635_, w_0838_, w_0640_);
not (w_0287_, w_0707_);
and (w_0314_, w_0405_, w_0494_);
and (w_0347_, in15[1], w_0474_);
and (w_0339_, w_0157_, w_0089_);
or (w_0731_, w_0686_, w_0619_);
and (w_0217_, w_0002_, w_0042_);
and (w_0117_, in15[0], w_0694_);
or (out10, w_0667_, w_0267_);
and (w_0444_, w_0598_, w_0680_);
and (w_0764_, w_0596_, w_0139_);
and (w_0150_, w_0554_, w_0434_);
and (w_0262_, in3[1], in4[0]);
or (w_0496_, in12[1], in11[1]);
and (w_0368_, w_0324_, w_0269_);
or (w_0471_, w_0155_, w_0111_);
or (w_0036_, w_0153_, w_0645_);
or (w_0558_, w_0307_, w_0437_);
or (w_0585_, w_0376_, w_0064_);
or (out1, w_0482_, w_0285_);
or (w_0140_, w_0274_, w_0319_);
and (w_0334_, w_0245_, w_0476_);
or (w_0189_, w_0443_, w_0310_);
or (w_0448_, w_0647_, w_0504_);
or (w_0233_, w_0581_, w_0503_);
and (w_0087_, w_0352_, w_0373_);
or (w_0335_, in15[0], w_0683_);
and (w_0793_, w_0202_, w_0514_);
and (w_0050_, w_0451_, w_0820_);
or (w_0209_, w_0546_, w_0146_);
or (w_0492_, w_0177_, w_0499_);
and (w_0499_, w_0351_, w_0234_);
and (w_0811_, w_0581_, w_0471_);
or (w_0425_, w_0166_, w_0586_);
and (w_0350_, w_0433_, w_0131_);
or (w_0545_, w_0026_, w_0792_);
or (w_0076_, w_0706_, w_0643_);
or (w_0049_, w_0577_, w_0676_);
and (w_0656_, w_0204_, w_0108_);
or (w_0509_, w_0604_, w_0145_);
and (w_0305_, in15[0], w_0207_);
not (w_0787_, in6[0]);
or (w_0020_, w_0355_, w_0278_);
or (w_0619_, w_0412_, w_0380_);
or (w_0240_, w_0800_, w_0245_);
or (w_0648_, w_0263_, w_0002_);
and (w_0232_, w_0054_, w_0529_);
or (w_0039_, w_0581_, w_0632_);
or (w_0841_, w_0063_, w_0787_);
or (w_0568_, w_0622_, w_0551_);
or (w_0293_, w_0568_, w_0298_);
and (w_0333_, w_0311_, w_0075_);
or (w_0820_, w_0440_, w_0790_);
and (w_0208_, w_0768_, w_0394_);
and (w_0657_, in1[1], in2[1]);
or (w_0717_, w_0046_, w_0738_);
and (w_0366_, w_0235_, w_0612_);
or (w_0164_, w_0003_, w_0107_);
and (w_0676_, w_0400_, w_0290_);
and (w_0647_, w_0712_, w_0228_);
and (w_0064_, w_0696_, w_0296_);
or (w_0061_, w_0054_, w_0529_);
or (w_0666_, w_0478_, w_0775_);
or (w_0344_, w_0120_, w_0378_);
or (w_0526_, w_0673_, w_0172_);
or (w_0342_, w_0235_, w_0612_);
or (w_0284_, w_0330_, w_0291_);
and (w_0521_, in11[0], in12[0]);
or (w_0612_, w_0569_, w_0769_);
or (w_0638_, w_0425_, w_0012_);
or (w_0436_, w_0215_, w_0133_);
or (w_0301_, w_0504_, w_0669_);
and (w_0336_, in5[0], in6[0]);
or (w_0707_, in14[1], in13[1]);
or (w_0354_, w_0203_, w_0596_);
and (w_0250_, in12[1], in11[1]);
or (w_0241_, w_0817_, w_0382_);
not (w_0476_, in11[1]);
and (w_0289_, in15[0], w_0547_);
or (w_0021_, w_0495_, w_0356_);
or (w_0723_, w_0672_, w_0458_);
or (w_0251_, w_0125_, w_0320_);
and (w_0198_, w_0598_, w_0363_);
or (w_0773_, w_0021_, w_0658_);
or (w_0300_, w_0215_, w_0441_);
or (w_0401_, w_0512_, w_0509_);
or (w_0292_, in15[0], w_0424_);
and (w_0621_, w_0180_, w_0237_);
not (w_0212_, w_0454_);
and (w_0329_, w_0781_, w_0099_);
or (w_0531_, w_0699_, w_0076_);
or (w_0119_, w_0510_, w_0344_);
and (w_0788_, w_0361_, w_0580_);
or (w_0306_, w_0677_, w_0796_);
or (w_0254_, w_0696_, w_0296_);
and (w_0817_, w_0191_, w_0201_);
and (w_0295_, w_0236_, w_0339_);
and (w_0431_, w_0345_, w_0331_);
or (w_0352_, w_0255_, w_0828_);
or (w_0007_, w_0295_, w_0465_);
and (w_0795_, w_0571_, w_0579_);
not (w_0631_, in1[0]);
and (w_0497_, w_0682_, w_0487_);
and (w_0291_, w_0096_, w_0735_);
not (w_0827_, in7[1]);
and (w_0572_, w_0504_, w_0506_);
or (w_0102_, in8[0], in7[1]);
not (w_0624_, w_0380_);
and (w_0740_, w_0227_, w_0196_);
and (w_0079_, w_0715_, w_0436_);
not (w_0770_, w_0809_);
and (w_0244_, in15[0], w_0635_);
and (w_0582_, w_0430_, w_0179_);
or (w_0761_, w_0047_, w_0741_);
and (w_0123_, in15[1], w_0527_);
and (w_0097_, w_0103_, w_0646_);
or (w_0091_, w_0581_, w_0471_);
and (w_0210_, w_0557_, w_0253_);
and (w_0744_, w_0240_, w_0236_);
and (w_0467_, w_0478_, w_0775_);
or (w_0227_, w_0255_, w_0338_);
and (w_0553_, w_0234_, w_0593_);
and (w_0109_, w_0568_, w_0707_);
and (w_0634_, w_0494_, w_0631_);
or (w_0194_, w_0445_, w_0407_);
or (w_0423_, w_0844_, w_0510_);
and (w_0312_, w_0132_, w_0822_);
or (w_0722_, w_0486_, w_0154_);
and (w_0361_, w_0054_, w_0457_);
and (w_0461_, w_0109_, w_0087_);
and (w_0383_, w_0080_, w_0122_);
or (w_0775_, w_0518_, w_0752_);
and (w_0759_, w_0496_, w_0415_);
not (w_0286_, w_0180_);
or (w_0668_, w_0582_, w_0650_);
and (w_0613_, w_0603_, w_0208_);
or (w_0345_, w_0581_, w_0085_);
or (w_0149_, in9[1], in10[0]);
and (w_0702_, w_0588_, w_0623_);
not (w_0766_, in6[1]);
or (w_0463_, w_0829_, w_0325_);
and (w_0591_, w_0732_, w_0463_);
or (w_0089_, w_0709_, w_0825_);
or (w_0828_, w_0477_, w_0795_);
or (w_0420_, in14[0], in13[1]);
and (w_0477_, w_0709_, w_0825_);
or (w_0832_, w_0720_, w_0040_);
not (w_0494_, in2[1]);
or (w_0270_, w_0581_, w_0241_);
and (w_0462_, w_0098_, w_0328_);
or (w_0328_, w_0305_, w_0753_);
or (w_0765_, w_0673_, w_0158_);
or (w_0729_, w_0080_, w_0515_);
and (w_0108_, w_0638_, w_0346_);
or (w_0593_, w_0737_, w_0748_);
not (w_0577_, w_0053_);
and (w_0282_, w_0370_, w_0674_);
and (w_0439_, w_0040_, w_0018_);
or (w_0721_, w_0500_, w_0303_);
and (w_0424_, w_0746_, w_0724_);
or (w_0712_, w_0361_, w_0580_);
or (w_0360_, w_0109_, w_0087_);
and (w_0672_, w_0452_, w_0109_);
and (w_0283_, w_0840_, w_0595_);
or (w_0324_, w_0281_, w_0084_);
not (w_0063_, in5[0]);
and (w_0317_, w_0797_, w_0116_);
or (w_0030_, w_0428_, w_0444_);
not (w_0750_, in14[0]);
and (w_0762_, w_0310_, w_0833_);
and (w_0814_, w_0406_, w_0206_);
or (w_0052_, w_0464_, w_0007_);
or (w_0570_, w_0141_, w_0446_);
not (w_0037_, w_0303_);
or (w_0512_, w_0334_, w_0250_);
or (w_0588_, w_0112_, w_0114_);
or (w_0413_, w_0812_, w_0478_);
or (w_0655_, w_0095_, w_0013_);
and (w_0470_, w_0734_, w_0153_);
or (w_0068_, w_0377_, w_0232_);
or (w_0121_, in9[1], in10[1]);
or (out7, w_0123_, w_0560_);
and (w_0330_, w_0799_, w_0780_);
and (w_0325_, w_0666_, w_0404_);
and (w_0501_, w_0581_, w_0074_);
or (w_0156_, w_0398_, w_0814_);
or (w_0288_, w_0314_, w_0657_);
and (w_0206_, w_0486_, w_0099_);
and (w_0017_, w_0407_, w_0151_);
and (w_0120_, w_0733_, w_0685_);
or (w_0603_, in13[0], in14[1]);
and (w_0205_, w_0250_, w_0280_);
and (w_0670_, w_0005_, w_0066_);
and (w_0308_, w_0570_, w_0379_);
or (w_0626_, w_0391_, w_0701_);
and (w_0154_, in3[1], in4[1]);
or (w_0434_, w_0121_, w_0742_);
or (w_0597_, w_0545_, w_0513_);
or (w_0105_, in15[0], w_0480_);
and (w_0363_, w_0197_, w_0428_);
or (w_0658_, w_0561_, w_0521_);
and (w_0725_, w_0348_, w_0797_);
and (w_0186_, w_0416_, w_0597_);
or (w_0661_, w_0159_, w_0743_);
not (w_0700_, w_0521_);
and (w_0567_, w_0161_, w_0591_);
and (w_0126_, w_0460_, w_0283_);
or (w_0812_, w_0516_, w_0537_);
or (w_0645_, w_0644_, w_0239_);
not (w_0066_, w_0198_);
or (w_0389_, in15[0], w_0137_);
or (out9, w_0628_, w_0642_);
and (w_0587_, w_0088_, w_0766_);
or (w_0428_, w_0653_, w_0166_);
and (w_0738_, w_0581_, w_0690_);
and (w_0479_, w_0313_, w_0512_);
or (w_0573_, w_0703_, w_0618_);
and (w_0692_, w_0415_, w_0636_);
and (w_0033_, w_0362_, w_0001_);
and (w_0048_, w_0836_, w_0627_);
or (w_0816_, w_0415_, w_0636_);
or (w_0124_, w_0126_, w_0534_);
not (w_0669_, w_0102_);
or (w_0633_, in15[0], w_0694_);
or (w_0754_, w_0149_, w_0397_);
and (w_0026_, w_0336_, w_0086_);
or (w_0054_, w_0405_, w_0815_);
and (w_0742_, w_0254_, w_0528_);
and (w_0022_, w_0098_, w_0442_);
or (w_0522_, w_0598_, w_0425_);
and (w_0706_, w_0571_, w_0535_);
and (w_0687_, w_0555_, w_0524_);
not (w_0800_, in11[0]);
and (w_0071_, w_0153_, w_0306_);
and (w_0453_, w_0119_, w_0384_);
or (w_0093_, w_0581_, w_0747_);
and (w_0225_, w_0765_, w_0727_);
or (w_0620_, w_0192_, w_0470_);
and (w_0104_, w_0049_, w_0386_);
or (w_0698_, in15[0], w_0635_);
or (w_0393_, in5[0], in6[0]);
not (w_0581_, in15[0]);
and (w_0168_, w_0264_, w_0520_);
and (w_0550_, w_0262_, w_0288_);
or (w_0734_, in7[1], in8[1]);
or (w_0682_, w_0425_, w_0444_);
and (w_0796_, w_0728_, w_0533_);
and (w_0772_, w_0033_, w_0081_);
and (w_0708_, w_0581_, w_0747_);
and (w_0417_, in7[0], in8[1]);
and (w_0340_, in15[1], w_0175_);
and (w_0058_, w_0581_, w_0124_);
or (w_0169_, w_0133_, w_0447_);
or (w_0566_, in15[0], w_0824_);
or (w_0486_, in1[0], in2[0]);
and (w_0195_, w_0512_, w_0509_);
and (w_0506_, w_0399_, w_0127_);
or (out4, w_0418_, w_0024_);
not (w_0435_, w_0136_);
and (w_0013_, w_0819_, w_0132_);
and (w_0515_, w_0818_, w_0072_);
and (w_0783_, w_0314_, w_0781_);
and (w_0159_, w_0720_, w_0185_);
and (w_0781_, in4[0], in3[0]);
not (w_0718_, w_0353_);
and (w_0265_, w_0307_, w_0437_);
or (w_0343_, w_0452_, w_0109_);
not (w_0405_, in1[1]);
and (w_0375_, w_0538_, w_0350_);
and (w_0737_, w_0274_, w_0804_);
and (w_0199_, w_0581_, w_0241_);
and (w_0556_, w_0215_, w_0832_);
or (out6, w_0808_, w_0789_);
and (w_0493_, w_0061_, w_0138_);
not (w_0245_, in12[1]);
or (w_0730_, w_0634_, w_0485_);
and (w_0319_, w_0688_, w_0751_);
or (w_0237_, in4[1], in3[0]);
or (w_0695_, w_0402_, w_0749_);
and (w_0495_, w_0468_, w_0829_);
or (w_0724_, w_0407_, w_0151_);
or (w_0178_, w_0728_, w_0301_);
and (w_0801_, w_0791_, w_0183_);
or (w_0010_, w_0250_, w_0280_);
and (w_0407_, w_0420_, w_0562_);
or (w_0798_, w_0571_, w_0353_);
and (w_0396_, w_0443_, w_0310_);
or (w_0652_, w_0318_, w_0490_);
and (w_0359_, w_0779_, w_0143_);
or (w_0507_, w_0641_, w_0240_);
or (w_0116_, w_0567_, w_0439_);
or (w_0132_, w_0715_, w_0417_);
and (w_0489_, w_0542_, w_0693_);
or (w_0822_, w_0656_, w_0760_);
and (w_0601_, w_0425_, w_0490_);
or (w_0555_, w_0271_, w_0803_);
or (w_0032_, w_0304_, w_0476_);
not (w_0561_, w_0171_);
and (w_0274_, w_0269_, w_0770_);
or (w_0118_, w_0654_, w_0725_);
and (w_0546_, in15[0], w_0491_);
or (w_0138_, w_0281_, w_0358_);
and (w_0719_, in15[0], w_0050_);
or (w_0277_, w_0469_, w_0090_);
or (w_0548_, w_0174_, w_0182_);
and (w_0808_, in15[1], w_0395_);
or (w_0782_, w_0779_, w_0143_);
or (w_0096_, w_0836_, w_0627_);
or (w_0697_, w_0589_, w_0275_);
and (w_0223_, w_0581_, w_0503_);
and (w_0518_, w_0274_, w_0319_);
and (w_0604_, w_0215_, w_0441_);
and (w_0753_, w_0581_, w_0723_);
or (w_0483_, w_0639_, w_0783_);
or (w_0171_, in11[0], in12[0]);
and (w_0008_, w_0055_, w_0607_);
or (w_0818_, w_0728_, w_0778_);
not (w_0586_, in3[0]);
and (w_0617_, w_0510_, w_0102_);
or (w_0711_, w_0581_, w_0690_);
or (w_0780_, w_0168_, w_0791_);
or (w_0429_, w_0316_, w_0176_);
not (w_0823_, in8[0]);
or (w_0674_, w_0336_, w_0086_);
and (w_0215_, in9[1], in10[0]);
or (w_0528_, w_0417_, w_0559_);
or (w_0456_, w_0658_, w_0541_);
or (w_0614_, w_0414_, w_0392_);
and (w_0769_, w_0112_, w_0114_);
or (w_0331_, in15[0], w_0590_);
or (w_0824_, w_0308_, w_0008_);
or (w_0777_, w_0679_, w_0615_);
or (w_0675_, w_0581_, w_0523_);
or (w_0170_, w_0262_, w_0288_);
and (w_0046_, in15[0], w_0381_);
and (w_0589_, in13[0], in14[1]);
or (w_0535_, w_0549_, w_0255_);
or (w_0520_, w_0733_, w_0721_);
or (w_0204_, in5[1], in6[1]);
or (w_0819_, w_0142_, w_0637_);
or (w_0290_, w_0180_, w_0237_);
and (w_0427_, in15[1], w_0793_);
and (w_0450_, w_0125_, w_0497_);
and (w_0465_, w_0255_, w_0828_);
and (w_0481_, w_0641_, w_0240_);
or (out3, w_0078_, w_0276_);
or (w_0768_, w_0313_, w_0512_);
and (w_0504_, in8[0], in7[1]);
or (w_0415_, w_0245_, w_0476_);
and (w_0683_, w_0806_, w_0354_);
or (w_0433_, w_0587_, w_0466_);
or (w_0732_, w_0051_, w_0574_);
and (w_0047_, w_0121_, w_0742_);
endmodule
