module new_sub_module1(
    input wire [2:0] new_in1,
    input wire [2:0] new_in2,
    input wire [2:0] new_in3,
    output wire [2:0] new_out1,
    output wire [2:0] new_out2
);
wire w_000_;
wire w_001_;
wire w_002_;
wire w_003_;
wire w_004_;
wire w_005_;
wire w_006_;
wire w_007_;
wire w_008_;
wire w_009_;
wire w_010_;
wire w_011_;
wire w_012_;
wire w_013_;
wire w_014_;
wire w_015_;
wire w_016_;
wire w_017_;
wire w_018_;
wire w_019_;
wire w_020_;
wire w_021_;
wire w_022_;
wire w_023_;
wire w_024_;
wire w_025_;
wire w_026_;
wire w_027_;
wire w_028_;
wire w_029_;
wire w_030_;
wire w_031_;
wire w_032_;
wire w_033_;
wire w_034_;
wire w_035_;
wire w_036_;
wire w_037_;
wire w_038_;
wire w_039_;
wire w_040_;
wire w_041_;
wire w_042_;
wire w_043_;
wire w_044_;
wire w_045_;
wire w_046_;
wire w_047_;
wire w_048_;
wire w_049_;
wire w_050_;
wire w_051_;
wire w_052_;
wire w_053_;
wire w_054_;
wire w_055_;
wire w_056_;
wire w_057_;
wire w_058_;
wire w_059_;
and (new_out2[0], w_001_, w_023_);
nand (w_055_, w_053_, w_016_);
nand (w_012_, w_008_, w_013_);
and (new_out1[0], w_029_, w_050_);
xor (w_054_, w_010_, w_006_);
and (w_037_, new_in1[1], w_049_);
and (w_020_, new_in1[1], new_in3[0]);
or (w_001_, w_018_, w_034_);
nand (w_009_, w_044_, w_036_);
xor (w_013_, new_in3[1], w_002_);
and (w_041_, new_in2[0], w_004_);
nand (w_034_, new_in2[2], w_053_);
and (w_030_, new_in3[2], new_in3[1]);
xor (w_043_, w_045_, w_015_);
xor (w_032_, w_020_, w_058_);
or (w_023_, w_053_, w_004_);
and (w_017_, new_in1[2], w_051_);
nand (w_014_, w_017_, w_038_);
xor (w_021_, w_031_, w_038_);
nor (w_042_, w_034_, w_011_);
not (w_025_, w_010_);
nand (w_039_, w_041_, w_059_);
not (w_022_, new_in2[0]);
nand (new_out2[1], w_024_, w_055_);
xor (w_010_, new_in2[0], new_in2[1]);
nand (w_007_, w_010_, w_048_);
or (w_036_, new_in3[1], w_008_);
nand (w_026_, w_025_, w_006_);
and (w_049_, new_in2[2], new_in3[2]);
not (w_051_, new_in3[1]);
xor (w_005_, w_028_, w_021_);
xor (w_035_, w_019_, w_054_);
and (w_011_, w_040_, w_000_);
or (w_057_, w_019_, w_054_);
xor (w_002_, w_041_, w_059_);
nand (w_044_, w_008_, w_002_);
nand (w_016_, w_012_, w_003_);
nand (new_out2[2], w_014_, w_033_);
and (w_015_, w_026_, w_057_);
and (w_003_, new_in2[2], w_027_);
and (new_out1[1], w_050_, w_035_);
and (w_000_, w_056_, w_009_);
nand (w_053_, new_in1[2], w_051_);
and (w_008_, new_in3[0], w_047_);
or (w_027_, w_008_, w_013_);
nor (w_019_, w_022_, new_in1[0]);
xor (w_048_, new_in1[1], w_049_);
xor (w_018_, new_in3[0], w_047_);
xor (w_029_, new_in2[0], new_in1[0]);
xor (w_038_, w_037_, w_030_);
and (w_028_, w_007_, w_039_);
nand (w_024_, w_017_, w_048_);
xor (w_058_, new_in1[2], new_in3[1]);
xor (w_040_, new_in3[2], w_005_);
nor (w_050_, new_in2[2], w_017_);
xor (w_045_, w_032_, w_031_);
xor (w_006_, new_in1[1], new_in3[0]);
and (w_046_, w_022_, new_in2[1]);
nand (w_056_, w_051_, w_002_);
and (w_004_, new_in1[1], new_in3[2]);
xor (w_059_, w_010_, w_048_);
and (new_out1[2], w_050_, w_043_);
xor (w_047_, new_in2[0], w_004_);
xor (w_031_, new_in2[2], w_046_);
nand (w_033_, w_052_, w_042_);
or (w_052_, w_040_, w_000_);
endmodule

module new_sub_module2(
    input wire [2:0] new_in1,
    input wire [2:0] new_in10,
    input wire [2:0] new_in11,
    input wire [2:0] new_in12,
    input wire [2:0] new_in2,
    input wire [2:0] new_in3,
    input wire [2:0] new_in4,
    input wire [2:0] new_in5,
    input wire [2:0] new_in6,
    input wire [2:0] new_in7,
    input wire [2:0] new_in8,
    input wire [2:0] new_in9,
    output wire [2:0] new_out1,
    output wire [2:0] new_out2,
    output wire [2:0] new_out3,
    output wire [2:0] new_out4,
    output wire [2:0] new_out5,
    output wire [2:0] new_out6
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
and (w_0444_, new_in6[0], new_in12[2]);
xor (w_0181_, w_0648_, w_0010_);
nand (w_0142_, w_0248_, w_0184_);
and (w_0390_, new_in4[2], new_in11[2]);
and (w_0460_, new_in5[0], new_in8[0]);
xor (w_0608_, w_0540_, w_0093_);
xor (w_0325_, w_0540_, w_0536_);
nand (w_0237_, w_0143_, w_0625_);
and (w_0248_, new_in7[0], new_in2[1]);
nand (w_0018_, w_0466_, w_0620_);
nand (w_0443_, w_0341_, w_0597_);
and (w_0165_, new_in5[1], new_in6[0]);
or (w_0104_, w_0036_, w_0576_);
or (w_0673_, w_0311_, w_0338_);
xor (w_0266_, w_0297_, w_0482_);
xor (w_0039_, new_in9[0], new_in3[0]);
and (w_0219_, w_0466_, w_0223_);
and (w_0117_, new_in5[0], new_in6[2]);
and (new_out4[1], w_0549_, w_0481_);
not (w_0100_, w_0329_);
not (w_0528_, new_in4[0]);
xor (w_0046_, new_in4[1], w_0360_);
nand (w_0340_, w_0391_, w_0361_);
xor (w_0586_, w_0392_, w_0413_);
nand (w_0365_, w_0323_, w_0102_);
and (w_0393_, new_in6[0], new_in1[0]);
xor (w_0145_, new_in6[1], w_0197_);
and (w_0624_, w_0435_, w_0120_);
nand (w_0008_, w_0423_, w_0642_);
and (w_0648_, w_0469_, w_0455_);
xor (w_0300_, w_0260_, w_0616_);
xor (w_0452_, w_0583_, w_0542_);
nand (w_0554_, new_in4[1], new_in2[1]);
and (w_0133_, w_0158_, w_0569_);
xor (w_0027_, new_in5[1], new_in8[1]);
nand (w_0280_, w_0427_, w_0007_);
nand (w_0307_, w_0383_, w_0644_);
xor (w_0234_, new_in5[0], w_0145_);
nand (w_0620_, w_0052_, w_0217_);
xor (w_0535_, w_0330_, w_0377_);
or (w_0435_, w_0478_, w_0315_);
xor (w_0063_, new_in9[2], w_0181_);
nand (w_0495_, new_in5[1], new_in10[1]);
and (w_0589_, w_0071_, w_0394_);
and (w_0583_, w_0165_, w_0646_);
nand (w_0077_, new_in6[1], new_in8[0]);
xor (w_0064_, w_0361_, w_0335_);
nand (w_0569_, w_0147_, w_0199_);
and (w_0184_, new_in7[1], new_in2[0]);
or (w_0594_, w_0367_, w_0275_);
xor (w_0590_, w_0650_, w_0214_);
and (w_0075_, new_in2[0], new_in4[0]);
and (w_0138_, w_0134_, w_0106_);
or (w_0004_, w_0190_, w_0564_);
xor (w_0475_, w_0375_, w_0091_);
and (w_0578_, w_0036_, w_0237_);
or (w_0440_, w_0036_, w_0233_);
xor (w_0558_, new_in10[2], w_0491_);
nand (w_0009_, new_in5[0], w_0491_);
nand (w_0038_, w_0021_, w_0205_);
nand (w_0344_, w_0036_, w_0112_);
and (w_0335_, new_in5[0], w_0294_);
xor (w_0168_, w_0503_, w_0590_);
and (w_0213_, w_0522_, w_0267_);
nand (w_0442_, w_0420_, w_0202_);
nand (w_0327_, new_in11[1], w_0026_);
or (w_0120_, w_0391_, w_0665_);
or (w_0132_, w_0036_, w_0446_);
xor (w_0458_, w_0049_, w_0250_);
and (w_0412_, w_0539_, w_0627_);
xor (w_0338_, w_0266_, w_0498_);
and (w_0062_, new_in5[0], w_0145_);
nand (w_0238_, w_0539_, w_0261_);
and (w_0424_, w_0438_, w_0580_);
or (w_0373_, w_0311_, w_0300_);
xor (w_0342_, new_in11[0], new_in4[0]);
xor (w_0033_, w_0107_, w_0332_);
and (w_0353_, w_0476_, w_0164_);
nand (w_0225_, w_0539_, w_0070_);
nand (w_0556_, w_0539_, w_0679_);
nand (w_0615_, w_0666_, w_0105_);
nand (w_0188_, w_0097_, w_0513_);
xor (w_0143_, new_in9[2], new_in10[2]);
or (w_0211_, w_0341_, w_0521_);
and (w_0140_, w_0466_, w_0176_);
or (w_0226_, w_0036_, w_0314_);
and (w_0593_, new_in12[0], new_in4[0]);
xor (w_0164_, new_in9[0], new_in10[0]);
and (w_0533_, w_0466_, w_0189_);
nand (w_0221_, w_0326_, w_0139_);
xor (w_0553_, w_0346_, w_0662_);
xor (w_0534_, w_0494_, w_0546_);
nand (w_0479_, w_0397_, w_0516_);
nand (w_0438_, w_0616_, w_0074_);
nand (w_0311_, new_in7[2], new_in2[0]);
xor (w_0262_, w_0177_, new_in2[2]);
nand (w_0497_, w_0143_, w_0328_);
and (w_0388_, w_0341_, w_0247_);
nand (w_0305_, w_0570_, w_0253_);
xor (w_0523_, new_in5[0], new_in10[0]);
and (new_out3[0], w_0645_, w_0065_);
and (w_0114_, w_0637_, w_0193_);
xor (w_0468_, new_in11[1], w_0026_);
xor (w_0343_, new_in11[2], w_0084_);
nand (w_0116_, w_0071_, w_0129_);
nand (w_0083_, w_0532_, w_0072_);
and (w_0392_, w_0068_, w_0426_);
xor (w_0048_, new_in5[1], new_in10[1]);
nand (w_0230_, new_in11[1], w_0285_);
nand (w_0163_, w_0353_, w_0033_);
nand (w_0663_, w_0259_, w_0320_);
or (w_0627_, w_0180_, w_0156_);
and (w_0021_, new_in9[2], new_in8[0]);
xor (w_0060_, w_0269_, w_0432_);
nand (w_0366_, w_0036_, w_0263_);
or (w_0426_, new_in1[2], new_in8[2]);
nand (w_0111_, w_0197_, w_0198_);
nand (w_0043_, new_in5[1], w_0286_);
xor (w_0001_, w_0446_, w_0207_);
xor (w_0260_, w_0555_, w_0155_);
nor (w_0476_, w_0385_, w_0293_);
xor (w_0135_, w_0588_, w_0628_);
nand (w_0095_, w_0246_, w_0148_);
nand (w_0414_, w_0036_, w_0527_);
xor (w_0603_, w_0135_, w_0076_);
or (w_0210_, w_0124_, w_0536_);
xor (w_0671_, w_0581_, new_in2[2]);
not (w_0581_, new_in7[1]);
xor (w_0324_, w_0049_, w_0622_);
nand (new_out3[2], w_0226_, w_0366_);
nand (w_0575_, w_0505_, w_0170_);
nand (w_0355_, w_0410_, w_0371_);
and (w_0137_, w_0389_, w_0080_);
nand (w_0264_, new_in1[2], w_0143_);
or (w_0445_, w_0094_, w_0047_);
xor (w_0400_, w_0585_, w_0517_);
nand (w_0112_, w_0264_, w_0019_);
nand (w_0115_, w_0367_, w_0396_);
nand (w_0000_, new_in9[1], new_in10[1]);
xor (w_0661_, w_0442_, w_0408_);
nand (w_0531_, w_0071_, w_0587_);
not (w_0297_, new_in11[0]);
nand (w_0525_, w_0058_, w_0005_);
xor (w_0073_, new_in12[0], w_0452_);
xor (w_0357_, new_in8[0], w_0310_);
xor (w_0488_, w_0292_, w_0553_);
and (w_0369_, w_0341_, w_0457_);
and (w_0377_, w_0607_, w_0083_);
or (w_0413_, w_0471_, w_0529_);
xor (w_0017_, new_in9[0], w_0471_);
nand (w_0515_, w_0573_, w_0412_);
xor (w_0592_, new_in9[1], w_0068_);
xor (w_0178_, w_0548_, w_0251_);
or (w_0341_, w_0476_, w_0107_);
or (w_0176_, w_0341_, w_0667_);
and (w_0124_, new_in7[0], w_0272_);
xor (w_0625_, new_in8[2], w_0275_);
and (w_0401_, w_0562_, w_0556_);
and (w_0222_, w_0407_, w_0465_);
xor (w_0349_, new_in9[0], new_in8[0]);
xor (w_0074_, w_0606_, w_0638_);
or (w_0612_, w_0434_, w_0090_);
and (w_0180_, new_in10[2], w_0491_);
nand (w_0602_, w_0341_, w_0305_);
nand (w_0196_, w_0071_, w_0362_);
xor (w_0322_, w_0528_, w_0456_);
nand (w_0035_, new_in11[2], w_0536_);
xor (w_0101_, w_0155_, w_0392_);
nand (w_0201_, w_0128_, w_0188_);
and (w_0119_, w_0319_, w_0490_);
xor (w_0619_, new_in4[1], new_in2[0]);
and (w_0579_, w_0539_, w_0514_);
and (w_0093_, new_in11[0], new_in4[0]);
xor (w_0191_, w_0290_, w_0108_);
xor (w_0198_, w_0391_, w_0361_);
nand (w_0622_, w_0030_, w_0510_);
xor (w_0477_, new_in10[1], new_in12[1]);
xor (w_0330_, w_0177_, w_0055_);
xor (w_0268_, new_in1[2], new_in6[2]);
nand (w_0637_, w_0231_, w_0507_);
nand (w_0483_, w_0551_, w_0545_);
nand (w_0641_, w_0522_, w_0552_);
xor (w_0621_, w_0167_, w_0592_);
and (w_0050_, new_in5[2], new_in12[0]);
nand (w_0319_, new_in6[1], w_0197_);
xor (w_0658_, new_in4[1], w_0362_);
and (w_0150_, w_0539_, w_0428_);
nand (w_0015_, w_0071_, w_0141_);
nand (w_0160_, w_0341_, w_0599_);
xor (w_0024_, w_0488_, w_0174_);
nor (w_0071_, w_0476_, w_0107_);
nand (w_0092_, w_0231_, w_0321_);
xor (w_0313_, w_0153_, w_0614_);
and (w_0241_, new_in6[1], new_in12[0]);
and (w_0303_, w_0382_, w_0249_);
nand (w_0012_, w_0143_, w_0651_);
nand (w_0146_, w_0143_, w_0454_);
nand (w_0203_, w_0309_, w_0633_);
nand (w_0500_, w_0423_, w_0099_);
nand (w_0068_, new_in1[2], new_in8[2]);
nand (w_0405_, w_0231_, w_0322_);
xor (w_0076_, w_0124_, w_0536_);
nand (w_0527_, w_0012_, w_0018_);
xor (w_0616_, w_0307_, w_0153_);
nand (w_0013_, new_in5[0], w_0286_);
xor (w_0517_, new_in8[1], new_in10[1]);
nand (w_0651_, w_0163_, w_0655_);
and (w_0385_, new_in1[0], new_in8[0]);
xor (w_0489_, w_0441_, w_0316_);
nand (w_0644_, w_0540_, w_0536_);
nand (w_0308_, w_0630_, w_0431_);
not (w_0418_, new_in11[1]);
nand (w_0229_, w_0341_, w_0429_);
nand (w_0374_, w_0116_, w_0409_);
xor (w_0482_, new_in6[0], new_in1[0]);
nand (w_0437_, w_0341_, w_0401_);
xor (w_0257_, new_in11[1], w_0285_);
xor (w_0010_, new_in5[2], new_in3[2]);
xor (w_0551_, new_in3[0], new_in12[0]);
xor (w_0040_, new_in7[2], w_0368_);
nand (w_0610_, w_0143_, w_0040_);
and (w_0269_, w_0606_, w_0638_);
xor (w_0380_, w_0029_, w_0145_);
and (w_0061_, w_0185_, w_0493_);
nand (w_0246_, w_0143_, w_0349_);
xor (w_0251_, w_0616_, w_0074_);
nand (w_0634_, w_0467_, w_0157_);
not (w_0296_, w_0045_);
nand (w_0306_, w_0311_, w_0641_);
nand (w_0081_, w_0273_, w_0160_);
xor (w_0587_, w_0525_, w_0337_);
xor (w_0314_, w_0195_, w_0136_);
xor (w_0668_, new_in5[2], new_in8[2]);
xor (w_0567_, w_0451_, w_0547_);
and (w_0228_, w_0238_, w_0560_);
xor (w_0281_, w_0248_, w_0184_);
xor (w_0187_, w_0397_, w_0516_);
nand (w_0570_, w_0231_, w_0676_);
xor (w_0016_, new_in5[1], w_0324_);
and (w_0529_, w_0385_, w_0107_);
nor (w_0107_, w_0471_, w_0113_);
xor (w_0110_, w_0222_, w_0268_);
nor (w_0113_, new_in1[1], new_in8[1]);
nand (w_0571_, w_0653_, w_0118_);
nand (new_out2[1], w_0243_, w_0082_);
xor (w_0653_, new_in7[0], new_in2[0]);
xor (w_0194_, w_0298_, w_0063_);
or (w_0645_, w_0036_, w_0001_);
nand (w_0420_, new_in10[1], new_in12[1]);
nand (w_0474_, w_0295_, w_0334_);
nand (w_0134_, w_0143_, w_0426_);
nand (w_0513_, w_0336_, w_0347_);
nand (w_0506_, w_0225_, w_0166_);
nand (w_0617_, w_0333_, w_0032_);
and (w_0309_, new_in8[0], w_0310_);
nand (w_0631_, w_0480_, w_0048_);
xor (w_0190_, w_0567_, w_0535_);
xor (w_0220_, w_0147_, w_0199_);
xor (w_0664_, w_0315_, w_0276_);
nand (w_0526_, w_0036_, w_0051_);
nand (w_0167_, new_in9[0], w_0471_);
nand (w_0079_, w_0232_, w_0257_);
xor (w_0546_, new_in11[1], new_in2[1]);
nand (w_0090_, w_0618_, w_0216_);
nand (w_0148_, w_0425_, w_0140_);
xor (w_0576_, w_0339_, w_0303_);
xor (w_0045_, new_in4[1], new_in11[1]);
nand (w_0271_, w_0341_, w_0114_);
and (new_out1[0], w_0103_, w_0254_);
xor (w_0066_, w_0475_, w_0137_);
xor (w_0434_, w_0309_, w_0633_);
and (w_0059_, new_in4[1], w_0362_);
xor (w_0439_, new_in12[2], new_in3[2]);
nand (w_0447_, new_in8[1], w_0270_);
xor (w_0153_, new_in7[2], new_in2[2]);
and (w_0473_, new_in11[0], w_0482_);
or (w_0623_, w_0304_, w_0520_);
xor (w_0411_, w_0278_, w_0299_);
xor (w_0337_, new_in7[2], new_in11[0]);
xor (w_0472_, new_in8[2], w_0194_);
xor (w_0277_, w_0241_, w_0057_);
and (new_out6[0], w_0089_, w_0132_);
and (w_0028_, w_0554_, w_0618_);
nand (w_0274_, w_0196_, w_0291_);
xor (w_0304_, w_0142_, w_0643_);
nand (w_0002_, new_in7[0], w_0143_);
nand (w_0067_, w_0486_, w_0574_);
nand (w_0591_, w_0231_, w_0621_);
nand (w_0502_, w_0577_, w_0283_);
or (w_0259_, w_0323_, w_0102_);
nand (w_0379_, w_0036_, w_0130_);
nand (w_0288_, w_0093_, w_0045_);
xor (w_0659_, w_0537_, w_0351_);
and (w_0240_, new_in4[1], w_0272_);
nand (w_0544_, w_0071_, w_0218_);
xor (w_0632_, new_in12[1], new_in3[1]);
xor (w_0368_, new_in8[0], new_in1[1]);
not (w_0278_, new_in5[1]);
and (w_0292_, w_0588_, w_0628_);
xor (w_0626_, w_0093_, w_0045_);
and (w_0352_, new_in7[0], new_in2[2]);
nand (w_0636_, w_0204_, w_0406_);
xor (w_0601_, w_0281_, w_0582_);
xor (w_0371_, new_in9[1], w_0598_);
xor (w_0250_, w_0622_, w_0439_);
nand (w_0618_, w_0075_, w_0519_);
or (w_0125_, w_0653_, w_0118_);
xor (w_0598_, w_0605_, w_0496_);
xor (w_0584_, w_0062_, w_0016_);
nand (w_0253_, w_0539_, w_0050_);
nand (w_0375_, w_0356_, w_0037_);
and (w_0094_, w_0266_, w_0498_);
xor (w_0541_, w_0181_, w_0208_);
nand (w_0639_, w_0511_, w_0602_);
nand (w_0563_, w_0473_, w_0468_);
and (w_0147_, new_in9[0], w_0523_);
nand (w_0295_, w_0539_, w_0182_);
nand (w_0394_, w_0304_, w_0520_);
xor (w_0536_, new_in7[1], new_in2[1]);
and (w_0320_, w_0231_, w_0365_);
nand (w_0103_, w_0126_, w_0404_);
not (w_0049_, new_in6[2]);
xor (w_0041_, w_0107_, w_0536_);
and (w_0367_, w_0009_, w_0395_);
nand (w_0097_, new_in9[1], new_in3[1]);
nand (new_out4[0], w_0008_, w_0200_);
xor (w_0290_, w_0551_, w_0545_);
and (w_0029_, new_in6[0], w_0551_);
or (w_0655_, w_0353_, w_0033_);
nand (w_0051_, w_0173_, w_0575_);
xor (w_0086_, w_0279_, w_0593_);
not (w_0294_, new_in6[0]);
xor (w_0347_, new_in9[1], new_in3[1]);
and (w_0227_, w_0660_, w_0258_);
nand (w_0036_, w_0566_, w_0151_);
nand (w_0263_, w_0596_, w_0610_);
nand (w_0356_, w_0418_, new_in2[1]);
nand (w_0600_, w_0539_, w_0239_);
xor (w_0224_, w_0397_, w_0664_);
nand (w_0429_, w_0673_, w_0056_);
xor (w_0323_, w_0472_, w_0096_);
nand (w_0158_, new_in9[1], w_0416_);
xor (w_0520_, w_0390_, w_0352_);
and (w_0149_, w_0503_, new_in10[2]);
xor (w_0055_, w_0572_, w_0668_);
xor (w_0561_, w_0476_, w_0653_);
and (w_0492_, w_0539_, w_0122_);
nand (new_out1[1], w_0500_, w_0414_);
xor (w_0456_, w_0467_, w_0157_);
nand (new_out5[1], w_0436_, w_0629_);
nand (w_0127_, new_in1[0], new_in8[0]);
xor (w_0635_, w_0023_, w_0444_);
xor (w_0464_, w_0240_, w_0403_);
xor (w_0354_, w_0143_, w_0392_);
nand (w_0298_, w_0317_, w_0355_);
nand (w_0398_, w_0460_, w_0027_);
nand (w_0183_, w_0539_, w_0236_);
nand (w_0058_, w_0177_, new_in2[1]);
and (w_0662_, w_0039_, w_0661_);
nand (w_0665_, w_0551_, w_0448_);
xor (w_0545_, new_in5[0], new_in6[0]);
nand (w_0524_, w_0071_, w_0608_);
nand (w_0599_, w_0006_, w_0255_);
xor (w_0091_, new_in11[2], new_in2[2]);
or (w_0499_, w_0036_, w_0584_);
nand (w_0372_, new_in5[1], new_in6[1]);
and (w_0614_, w_0035_, w_0634_);
xor (w_0208_, w_0453_, w_0635_);
xor (w_0559_, w_0380_, w_0220_);
xor (w_0159_, new_in8[1], w_0164_);
and (w_0205_, new_in7[0], new_in12[0]);
and (w_0652_, w_0230_, w_0079_);
or (w_0189_, w_0341_, w_0658_);
xor (w_0026_, w_0393_, w_0557_);
nand (w_0179_, w_0231_, w_0017_);
xor (w_0315_, w_0165_, w_0646_);
xor (w_0370_, w_0109_, w_0384_);
and (w_0611_, w_0433_, w_0479_);
nand (w_0105_, w_0466_, w_0422_);
and (w_0654_, new_in9[0], new_in10[0]);
nand (w_0247_, w_0127_, w_0231_);
or (w_0042_, w_0290_, w_0036_);
not (w_0209_, new_in6[1]);
xor (w_0656_, w_0060_, w_0424_);
xor (w_0496_, new_in5[1], new_in3[1]);
xor (w_0129_, w_0059_, w_0011_);
nand (w_0649_, w_0036_, w_0615_);
nand (w_0465_, w_0393_, w_0557_);
not (w_0478_, w_0197_);
nand (w_0151_, w_0430_, w_0624_);
nand (w_0511_, w_0071_, w_0066_);
and (w_0678_, new_in11[2], new_in4[0]);
xor (w_0072_, new_in4[1], w_0613_);
or (w_0674_, w_0341_, w_0601_);
xor (w_0677_, w_0152_, w_0169_);
not (w_0162_, w_0476_);
nand (w_0514_, w_0190_, w_0564_);
or (w_0122_, w_0164_, w_0367_);
xor (w_0461_, w_0651_, w_0659_);
nand (w_0255_, w_0004_, w_0579_);
or (w_0005_, w_0240_, w_0403_);
nand (w_0383_, new_in7[1], new_in2[1]);
nand (w_0014_, w_0470_, w_0373_);
nand (w_0574_, w_0143_, w_0672_);
nand (w_0486_, w_0466_, w_0374_);
and (w_0480_, new_in5[0], new_in10[0]);
nand (w_0530_, w_0539_, w_0154_);
nand (w_0032_, w_0271_, w_0219_);
and (w_0467_, new_in11[1], w_0653_);
xor (w_0136_, w_0168_, w_0133_);
xor (w_0359_, w_0113_, w_0000_);
nand (w_0056_, w_0311_, w_0284_);
and (w_0628_, w_0039_, w_0258_);
and (w_0504_, new_in9[1], new_in6[2]);
xor (w_0408_, new_in10[2], new_in12[2]);
and (w_0351_, w_0025_, w_0163_);
or (w_0675_, w_0311_, w_0558_);
nand (w_0490_, w_0029_, w_0145_);
and (w_0395_, w_0043_, w_0034_);
xor (w_0258_, w_0088_, w_0477_);
nand (w_0019_, w_0466_, w_0081_);
xor (w_0633_, new_in8[1], w_0270_);
not (w_0423_, w_0036_);
nand (w_0331_, w_0231_, w_0487_);
and (w_0532_, new_in4[0], w_0078_);
not (w_0503_, new_in9[2]);
nand (w_0089_, w_0502_, w_0485_);
or (w_0321_, new_in11[1], w_0653_);
nand (w_0080_, w_0059_, w_0011_);
nand (w_0564_, w_0020_, w_0445_);
nand (w_0333_, w_0143_, w_0359_);
or (w_0609_, w_0467_, w_0092_);
or (w_0245_, w_0367_, w_0595_);
xor (w_0487_, w_0342_, w_0561_);
nand (w_0431_, w_0466_, w_0235_);
and (w_0572_, w_0302_, w_0398_);
nor (w_0293_, new_in1[0], new_in8[0]);
nand (w_0505_, w_0341_, w_0192_);
xor (w_0197_, w_0312_, w_0632_);
xor (w_0155_, new_in4[2], new_in11[2]);
or (w_0252_, w_0626_, w_0325_);
or (w_0436_, w_0036_, w_0191_);
nand (w_0406_, w_0466_, w_0123_);
not (w_0242_, new_in10[0]);
nand (w_0131_, w_0036_, w_0350_);
xor (w_0085_, w_0272_, new_in4[0]);
xor (w_0521_, w_0093_, w_0325_);
nand (w_0212_, w_0372_, w_0340_);
and (w_0360_, new_in4[0], w_0456_);
and (w_0547_, w_0327_, w_0563_);
xor (w_0403_, new_in4[2], new_in2[1]);
nand (w_0463_, w_0450_, w_0533_);
xor (w_0047_, w_0161_, w_0329_);
nand (w_0350_, w_0264_, w_0287_);
xor (w_0169_, new_in5[2], new_in6[2]);
nand (w_0317_, new_in9[1], w_0598_);
xor (w_0310_, new_in9[0], w_0441_);
nand (new_out3[1], w_0415_, w_0175_);
nand (w_0409_, w_0647_, w_0417_);
and (w_0282_, w_0466_, w_0531_);
or (w_0223_, w_0341_, w_0464_);
and (w_0057_, new_in6[0], new_in12[1]);
xor (w_0141_, w_0304_, w_0260_);
xor (w_0199_, new_in9[1], w_0416_);
xor (w_0270_, w_0410_, w_0371_);
nand (w_0629_, w_0036_, w_0095_);
and (w_0585_, new_in9[0], new_in8[0]);
xor (w_0660_, w_0336_, w_0347_);
xor (w_0174_, w_0153_, w_0501_);
xor (w_0640_, w_0611_, w_0073_);
or (w_0031_, w_0341_, w_0178_);
xor (w_0396_, w_0127_, w_0107_);
nand (w_0381_, w_0036_, w_0138_);
and (w_0605_, new_in5[0], new_in3[0]);
nand (w_0289_, w_0036_, w_0308_);
nand (w_0670_, w_0550_, w_0492_);
xor (w_0161_, w_0473_, w_0468_);
or (w_0326_, w_0341_, w_0619_);
nand (w_0152_, w_0376_, w_0265_);
nand (w_0453_, w_0241_, w_0057_);
xor (w_0613_, w_0460_, w_0027_);
nand (w_0144_, w_0423_, w_0234_);
nand (w_0647_, w_0231_, w_0069_);
xor (w_0595_, w_0143_, w_0206_);
and (w_0391_, new_in5[0], new_in6[0]);
nand (w_0428_, w_0626_, w_0325_);
nand (new_out5[0], w_0042_, w_0131_);
or (w_0348_, w_0036_, w_0541_);
xor (w_0108_, w_0197_, w_0064_);
nand (w_0030_, new_in12[1], new_in3[1]);
and (w_0606_, new_in4[1], new_in11[0]);
nand (w_0364_, w_0231_, w_0603_);
xor (w_0557_, new_in6[1], new_in1[1]);
nand (w_0382_, w_0315_, w_0276_);
and (w_0646_, new_in5[0], new_in6[1]);
nand (w_0192_, w_0405_, w_0530_);
nand (w_0560_, w_0483_, w_0231_);
and (w_0650_, w_0495_, w_0631_);
not (w_0177_, new_in4[2]);
and (w_0299_, new_in6[2], w_0538_);
xor (w_0256_, new_in9[1], new_in10[1]);
xor (w_0432_, w_0582_, w_0678_);
and (w_0232_, new_in11[0], new_in2[0]);
nand (w_0204_, w_0143_, w_0159_);
nand (w_0358_, w_0071_, w_0172_);
xor (w_0421_, w_0038_, w_0086_);
nand (w_0596_, w_0466_, w_0639_);
xor (w_0102_, w_0028_, w_0262_);
nand (w_0287_, w_0466_, w_0186_);
nand (w_0481_, w_0044_, w_0578_);
nand (w_0023_, new_in6[1], new_in12[1]);
xor (w_0157_, new_in11[2], w_0536_);
xor (w_0328_, w_0293_, w_0654_);
and (w_0007_, w_0036_, w_0466_);
nand (w_0607_, new_in4[1], w_0613_);
and (w_0170_, w_0466_, w_0031_);
xor (w_0509_, w_0169_, w_0212_);
or (w_0449_, w_0290_, w_0108_);
nor (w_0054_, w_0483_, w_0111_);
nand (w_0053_, w_0654_, w_0256_);
nand (new_out5[2], w_0440_, w_0289_);
nand (w_0577_, w_0670_, w_0301_);
xor (w_0672_, new_in7[1], new_in1[0]);
or (w_0549_, w_0036_, w_0224_);
xor (w_0084_, w_0248_, w_0671_);
nand (w_0457_, w_0539_, w_0504_);
nand (w_0470_, w_0231_, w_0370_);
nand (w_0669_, w_0612_, w_0213_);
xor (w_0195_, w_0119_, w_0458_);
xor (w_0172_, w_0343_, w_0652_);
not (w_0272_, new_in2[0]);
nand (new_out6[2], w_0499_, w_0280_);
and (w_0638_, new_in11[1], new_in4[0]);
nand (w_0186_, w_0544_, w_0378_);
xor (w_0218_, w_0540_, w_0342_);
xor (w_0099_, w_0598_, w_0277_);
nand (w_0407_, new_in6[1], new_in1[1]);
nand (w_0484_, w_0341_, w_0014_);
nand (w_0154_, w_0115_, w_0594_);
xor (w_0275_, w_0654_, w_0256_);
nand (new_out1[2], w_0348_, w_0649_);
and (w_0410_, new_in9[0], w_0441_);
xor (w_0332_, w_0256_, w_0657_);
xor (w_0128_, new_in10[0], new_in12[0]);
xor (w_0069_, w_0296_, w_0041_);
and (w_0096_, w_0447_, w_0203_);
xor (w_0261_, w_0342_, w_0653_);
xor (w_0339_, w_0452_, w_0508_);
and (new_out2[2], w_0381_, w_0512_);
nand (w_0459_, w_0087_, w_0663_);
nand (w_0249_, w_0397_, w_0664_);
nand (w_0450_, w_0331_, w_0369_);
nand (w_0193_, w_0252_, w_0150_);
nand (w_0020_, w_0161_, w_0100_);
nand (w_0402_, w_0013_, w_0573_);
nand (w_0267_, w_0434_, w_0090_);
nand (w_0493_, w_0171_, new_in10[1]);
nand (w_0025_, w_0107_, w_0332_);
nand (w_0052_, w_0071_, w_0244_);
nand (new_out6[1], w_0144_, w_0526_);
nand (w_0419_, w_0367_, w_0586_);
and (w_0283_, w_0466_, w_0211_);
nand (w_0550_, w_0162_, w_0367_);
and (w_0236_, new_in8[0], new_in12[0]);
nand (w_0006_, w_0231_, w_0024_);
nand (w_0202_, w_0088_, w_0477_);
and (w_0399_, w_0539_, w_0363_);
or (w_0216_, w_0075_, w_0519_);
xor (w_0508_, new_in12[1], w_0565_);
nand (w_0573_, w_0180_, w_0156_);
nand (w_0666_, w_0143_, w_0461_);
xor (w_0543_, w_0313_, w_0046_);
xor (w_0542_, w_0372_, w_0117_);
xor (w_0643_, w_0539_, w_0383_);
xor (w_0182_, w_0402_, w_0411_);
xor (w_0667_, w_0281_, w_0626_);
or (w_0376_, w_0361_, w_0335_);
and (w_0491_, new_in6[0], w_0312_);
nand (w_0243_, w_0423_, w_0187_);
xor (w_0207_, new_in9[0], w_0523_);
nand (w_0217_, w_0341_, w_0506_);
nand (w_0430_, w_0452_, w_0250_);
xor (w_0070_, w_0021_, w_0205_);
nand (w_0173_, new_in9[1], w_0149_);
nand (w_0175_, w_0036_, w_0067_);
xor (w_0329_, w_0532_, w_0072_);
nand (w_0318_, w_0071_, w_0656_);
nand (w_0389_, new_in4[2], w_0534_);
and (w_0098_, w_0522_, w_0571_);
nand (w_0510_, w_0312_, w_0632_);
nand (w_0265_, w_0278_, new_in6[1]);
nand (w_0630_, w_0143_, w_0400_);
and (w_0404_, w_0036_, w_0146_);
or (w_0254_, w_0036_, w_0489_);
nand (w_0582_, new_in4[1], new_in11[1]);
and (w_0334_, w_0341_, w_0591_);
nand (w_0422_, w_0358_, w_0387_);
and (w_0485_, w_0036_, w_0345_);
nor (w_0286_, w_0209_, w_0030_);
xor (w_0346_, w_0201_, w_0227_);
xor (w_0276_, new_in12[0], new_in3[2]);
and (w_0206_, w_0000_, w_0053_);
and (w_0548_, w_0093_, w_0325_);
or (w_0037_, w_0494_, w_0546_);
and (w_0417_, w_0341_, w_0600_);
or (w_0507_, w_0054_, w_0109_);
nand (w_0469_, new_in5[1], new_in3[1]);
xor (w_0552_, w_0357_, w_0085_);
nand (w_0562_, w_0231_, w_0543_);
xor (w_0462_, w_0250_, w_0677_);
and (w_0215_, w_0463_, w_0002_);
xor (w_0233_, w_0449_, w_0462_);
xor (w_0285_, new_in7[0], new_in2[1]);
nand (w_0044_, w_0466_, w_0022_);
nand (w_0106_, w_0484_, w_0282_);
xor (w_0446_, new_in6[0], w_0551_);
nand (new_out4[2], w_0104_, w_0344_);
and (w_0312_, new_in3[0], new_in12[0]);
nand (w_0139_, w_0341_, w_0228_);
xor (w_0516_, new_in3[2], w_0315_);
and (w_0121_, new_in7[0], new_in9[2]);
and (w_0539_, new_in7[2], new_in2[0]);
xor (w_0361_, new_in5[1], new_in6[1]);
nand (w_0501_, w_0518_, w_0210_);
nand (new_out2[0], w_0008_, w_0379_);
nand (w_0433_, new_in3[2], w_0315_);
or (w_0512_, w_0036_, w_0640_);
or (w_0566_, w_0452_, w_0250_);
nand (w_0387_, w_0341_, w_0459_);
nand (w_0022_, w_0674_, w_0443_);
nand (w_0455_, w_0605_, w_0496_);
nand (w_0034_, new_in5[2], w_0299_);
and (w_0301_, w_0341_, w_0609_);
nand (w_0239_, new_in3[0], new_in10[0]);
nand (w_0273_, w_0623_, w_0589_);
not (w_0171_, new_in9[1]);
and (w_0397_, new_in3[1], w_0391_);
nand (w_0166_, w_0311_, w_0669_);
and (w_0130_, w_0003_, w_0497_);
nand (w_0604_, w_0183_, w_0306_);
and (w_0540_, new_in7[0], new_in2[0]);
nand (w_0425_, w_0515_, w_0568_);
xor (w_0078_, new_in5[0], new_in8[0]);
nand (w_0123_, w_0524_, w_0229_);
nand (w_0345_, w_0143_, w_0392_);
xor (w_0244_, w_0232_, w_0257_);
nand (w_0200_, w_0036_, w_0636_);
xor (w_0011_, new_in4[2], w_0534_);
xor (w_0642_, new_in3[1], w_0391_);
nand (w_0378_, w_0675_, w_0388_);
and (w_0494_, new_in11[0], w_0272_);
nand (w_0518_, w_0581_, new_in2[1]);
nand (w_0427_, w_0318_, w_0437_);
and (w_0088_, new_in10[0], new_in12[0]);
xor (w_0362_, new_in11[0], new_in2[0]);
nand (w_0580_, w_0548_, w_0251_);
nand (w_0555_, w_0582_, w_0288_);
nand (w_0363_, w_0094_, w_0047_);
or (w_0522_, new_in4[2], new_in11[2]);
and (w_0679_, w_0245_, w_0419_);
and (w_0231_, w_0311_, w_0522_);
and (w_0657_, new_in9[0], w_0242_);
nand (w_0284_, w_0125_, w_0098_);
nand (w_0597_, w_0364_, w_0386_);
nand (w_0415_, w_0423_, w_0559_);
nand (w_0087_, w_0539_, w_0421_);
xor (w_0537_, w_0061_, w_0354_);
and (w_0471_, new_in1[1], new_in8[1]);
xor (w_0416_, w_0480_, w_0048_);
and (w_0538_, new_in12[2], new_in3[2]);
and (w_0109_, w_0483_, w_0111_);
nand (w_0386_, w_0445_, w_0399_);
xor (w_0676_, w_0153_, w_0101_);
and (w_0568_, w_0341_, w_0179_);
and (w_0588_, w_0128_, w_0660_);
xor (w_0451_, new_in11[2], w_0110_);
nand (w_0003_, w_0466_, w_0221_);
xor (w_0498_, new_in4[0], w_0078_);
not (w_0466_, w_0143_);
nand (w_0118_, w_0128_, w_0039_);
and (w_0336_, new_in9[0], new_in3[0]);
nand (w_0082_, w_0036_, w_0617_);
or (w_0185_, w_0256_, w_0657_);
xor (w_0441_, new_in5[0], new_in3[0]);
nand (w_0302_, new_in5[1], new_in8[1]);
nand (w_0291_, w_0341_, w_0604_);
nand (w_0565_, new_in12[0], new_in3[2]);
nand (w_0065_, w_0036_, w_0215_);
xor (w_0519_, new_in4[1], new_in2[1]);
xor (w_0156_, new_in5[0], w_0286_);
nand (w_0448_, w_0478_, w_0315_);
and (w_0384_, w_0250_, w_0509_);
xor (w_0279_, w_0077_, w_0121_);
and (w_0316_, new_in6[0], new_in12[0]);
xor (w_0214_, new_in5[2], new_in10[2]);
nand (w_0235_, w_0015_, w_0474_);
nand (w_0126_, w_0466_, w_0274_);
xor (w_0454_, w_0476_, w_0164_);
endmodule

module new_sub_module3(
    input wire [1:0] new_in11,
    input wire [1:0] new_in7,
    input wire [6:0] new_in1,
    input wire [6:0] new_in10,
    input wire [6:0] new_in3,
    input wire [6:0] new_in8,
    input wire [6:0] new_in9,
    input wire [8:0] new_in2,
    input wire [8:0] new_in4,
    input wire [8:0] new_in5,
    input wire [8:0] new_in6,
    output wire [3:0] new_out1,
    output wire [3:0] new_out10,
    output wire [3:0] new_out11,
    output wire [3:0] new_out3,
    output wire [3:0] new_out5,
    output wire [3:0] new_out6,
    output wire [3:0] new_out7,
    output wire [3:0] new_out8,
    output wire [3:0] new_out9,
    output wire new_out2,
    output wire new_out4
);
wire w_0000_;
wire w_0001_;
wire w_0002_;
wire w_0003_;
wire w_0004_;
wire w_0005_;
wire w_0006_;
wire w_0007_;
wire w_0008_;
wire w_0009_;
wire w_0010_;
wire w_0011_;
wire w_0012_;
wire w_0013_;
wire w_0014_;
wire w_0015_;
wire w_0016_;
wire w_0017_;
wire w_0018_;
wire w_0019_;
wire w_0020_;
wire w_0021_;
wire w_0022_;
wire w_0023_;
wire w_0024_;
wire w_0025_;
wire w_0026_;
wire w_0027_;
wire w_0028_;
wire w_0029_;
wire w_0030_;
wire w_0031_;
wire w_0032_;
wire w_0033_;
wire w_0034_;
wire w_0035_;
wire w_0036_;
wire w_0037_;
wire w_0038_;
wire w_0039_;
wire w_0040_;
wire w_0041_;
wire w_0042_;
wire w_0043_;
wire w_0044_;
wire w_0045_;
wire w_0046_;
wire w_0047_;
wire w_0048_;
wire w_0049_;
wire w_0050_;
wire w_0051_;
wire w_0052_;
wire w_0053_;
wire w_0054_;
wire w_0055_;
wire w_0056_;
wire w_0057_;
wire w_0058_;
wire w_0059_;
wire w_0060_;
wire w_0061_;
wire w_0062_;
wire w_0063_;
wire w_0064_;
wire w_0065_;
wire w_0066_;
wire w_0067_;
wire w_0068_;
wire w_0069_;
wire w_0070_;
wire w_0071_;
wire w_0072_;
wire w_0073_;
wire w_0074_;
wire w_0075_;
wire w_0076_;
wire w_0077_;
wire w_0078_;
wire w_0079_;
wire w_0080_;
wire w_0081_;
wire w_0082_;
wire w_0083_;
wire w_0084_;
wire w_0085_;
wire w_0086_;
wire w_0087_;
wire w_0088_;
wire w_0089_;
wire w_0090_;
wire w_0091_;
wire w_0092_;
wire w_0093_;
wire w_0094_;
wire w_0095_;
wire w_0096_;
wire w_0097_;
wire w_0098_;
wire w_0099_;
wire w_0100_;
wire w_0101_;
wire w_0102_;
wire w_0103_;
wire w_0104_;
wire w_0105_;
wire w_0106_;
wire w_0107_;
wire w_0108_;
wire w_0109_;
wire w_0110_;
wire w_0111_;
wire w_0112_;
wire w_0113_;
wire w_0114_;
wire w_0115_;
wire w_0116_;
wire w_0117_;
wire w_0118_;
wire w_0119_;
wire w_0120_;
wire w_0121_;
wire w_0122_;
wire w_0123_;
wire w_0124_;
wire w_0125_;
wire w_0126_;
wire w_0127_;
wire w_0128_;
wire w_0129_;
wire w_0130_;
wire w_0131_;
wire w_0132_;
wire w_0133_;
wire w_0134_;
wire w_0135_;
wire w_0136_;
wire w_0137_;
wire w_0138_;
wire w_0139_;
wire w_0140_;
wire w_0141_;
wire w_0142_;
wire w_0143_;
wire w_0144_;
wire w_0145_;
wire w_0146_;
wire w_0147_;
wire w_0148_;
wire w_0149_;
wire w_0150_;
wire w_0151_;
wire w_0152_;
wire w_0153_;
wire w_0154_;
wire w_0155_;
wire w_0156_;
wire w_0157_;
wire w_0158_;
wire w_0159_;
wire w_0160_;
wire w_0161_;
wire w_0162_;
wire w_0163_;
wire w_0164_;
wire w_0165_;
wire w_0166_;
wire w_0167_;
wire w_0168_;
wire w_0169_;
wire w_0170_;
wire w_0171_;
wire w_0172_;
wire w_0173_;
wire w_0174_;
wire w_0175_;
wire w_0176_;
wire w_0177_;
wire w_0178_;
wire w_0179_;
wire w_0180_;
wire w_0181_;
wire w_0182_;
wire w_0183_;
wire w_0184_;
wire w_0185_;
wire w_0186_;
wire w_0187_;
wire w_0188_;
wire w_0189_;
wire w_0190_;
wire w_0191_;
wire w_0192_;
wire w_0193_;
wire w_0194_;
wire w_0195_;
wire w_0196_;
wire w_0197_;
wire w_0198_;
wire w_0199_;
wire w_0200_;
wire w_0201_;
wire w_0202_;
wire w_0203_;
wire w_0204_;
wire w_0205_;
wire w_0206_;
wire w_0207_;
wire w_0208_;
wire w_0209_;
wire w_0210_;
wire w_0211_;
wire w_0212_;
wire w_0213_;
wire w_0214_;
wire w_0215_;
wire w_0216_;
wire w_0217_;
wire w_0218_;
wire w_0219_;
wire w_0220_;
wire w_0221_;
wire w_0222_;
wire w_0223_;
wire w_0224_;
wire w_0225_;
wire w_0226_;
wire w_0227_;
wire w_0228_;
wire w_0229_;
wire w_0230_;
wire w_0231_;
wire w_0232_;
wire w_0233_;
wire w_0234_;
wire w_0235_;
wire w_0236_;
wire w_0237_;
wire w_0238_;
wire w_0239_;
wire w_0240_;
wire w_0241_;
wire w_0242_;
wire w_0243_;
wire w_0244_;
wire w_0245_;
wire w_0246_;
wire w_0247_;
wire w_0248_;
wire w_0249_;
wire w_0250_;
wire w_0251_;
wire w_0252_;
wire w_0253_;
wire w_0254_;
wire w_0255_;
wire w_0256_;
wire w_0257_;
wire w_0258_;
wire w_0259_;
wire w_0260_;
wire w_0261_;
wire w_0262_;
wire w_0263_;
wire w_0264_;
wire w_0265_;
wire w_0266_;
wire w_0267_;
wire w_0268_;
wire w_0269_;
wire w_0270_;
wire w_0271_;
wire w_0272_;
wire w_0273_;
wire w_0274_;
wire w_0275_;
wire w_0276_;
wire w_0277_;
wire w_0278_;
wire w_0279_;
wire w_0280_;
wire w_0281_;
wire w_0282_;
wire w_0283_;
wire w_0284_;
wire w_0285_;
wire w_0286_;
wire w_0287_;
wire w_0288_;
wire w_0289_;
wire w_0290_;
wire w_0291_;
wire w_0292_;
wire w_0293_;
wire w_0294_;
wire w_0295_;
wire w_0296_;
wire w_0297_;
wire w_0298_;
wire w_0299_;
wire w_0300_;
wire w_0301_;
wire w_0302_;
wire w_0303_;
wire w_0304_;
wire w_0305_;
wire w_0306_;
wire w_0307_;
wire w_0308_;
wire w_0309_;
wire w_0310_;
wire w_0311_;
wire w_0312_;
wire w_0313_;
wire w_0314_;
wire w_0315_;
wire w_0316_;
wire w_0317_;
wire w_0318_;
wire w_0319_;
wire w_0320_;
wire w_0321_;
wire w_0322_;
wire w_0323_;
wire w_0324_;
wire w_0325_;
wire w_0326_;
wire w_0327_;
wire w_0328_;
wire w_0329_;
wire w_0330_;
wire w_0331_;
wire w_0332_;
wire w_0333_;
wire w_0334_;
wire w_0335_;
wire w_0336_;
wire w_0337_;
wire w_0338_;
wire w_0339_;
wire w_0340_;
wire w_0341_;
wire w_0342_;
wire w_0343_;
wire w_0344_;
wire w_0345_;
wire w_0346_;
wire w_0347_;
wire w_0348_;
wire w_0349_;
wire w_0350_;
wire w_0351_;
wire w_0352_;
wire w_0353_;
wire w_0354_;
wire w_0355_;
wire w_0356_;
wire w_0357_;
wire w_0358_;
wire w_0359_;
wire w_0360_;
wire w_0361_;
wire w_0362_;
wire w_0363_;
wire w_0364_;
wire w_0365_;
wire w_0366_;
wire w_0367_;
wire w_0368_;
wire w_0369_;
wire w_0370_;
wire w_0371_;
wire w_0372_;
wire w_0373_;
wire w_0374_;
wire w_0375_;
wire w_0376_;
wire w_0377_;
wire w_0378_;
wire w_0379_;
wire w_0380_;
wire w_0381_;
wire w_0382_;
wire w_0383_;
wire w_0384_;
wire w_0385_;
wire w_0386_;
wire w_0387_;
wire w_0388_;
wire w_0389_;
wire w_0390_;
wire w_0391_;
wire w_0392_;
wire w_0393_;
wire w_0394_;
wire w_0395_;
wire w_0396_;
wire w_0397_;
wire w_0398_;
wire w_0399_;
wire w_0400_;
wire w_0401_;
wire w_0402_;
wire w_0403_;
wire w_0404_;
wire w_0405_;
wire w_0406_;
wire w_0407_;
wire w_0408_;
wire w_0409_;
wire w_0410_;
wire w_0411_;
wire w_0412_;
wire w_0413_;
wire w_0414_;
wire w_0415_;
wire w_0416_;
wire w_0417_;
wire w_0418_;
wire w_0419_;
wire w_0420_;
wire w_0421_;
wire w_0422_;
wire w_0423_;
wire w_0424_;
wire w_0425_;
wire w_0426_;
wire w_0427_;
wire w_0428_;
wire w_0429_;
wire w_0430_;
wire w_0431_;
wire w_0432_;
wire w_0433_;
wire w_0434_;
wire w_0435_;
wire w_0436_;
wire w_0437_;
wire w_0438_;
wire w_0439_;
wire w_0440_;
wire w_0441_;
wire w_0442_;
wire w_0443_;
wire w_0444_;
wire w_0445_;
wire w_0446_;
wire w_0447_;
wire w_0448_;
wire w_0449_;
wire w_0450_;
wire w_0451_;
wire w_0452_;
wire w_0453_;
wire w_0454_;
wire w_0455_;
wire w_0456_;
wire w_0457_;
wire w_0458_;
wire w_0459_;
wire w_0460_;
wire w_0461_;
wire w_0462_;
wire w_0463_;
wire w_0464_;
wire w_0465_;
wire w_0466_;
wire w_0467_;
wire w_0468_;
wire w_0469_;
wire w_0470_;
wire w_0471_;
wire w_0472_;
wire w_0473_;
wire w_0474_;
wire w_0475_;
wire w_0476_;
wire w_0477_;
wire w_0478_;
wire w_0479_;
wire w_0480_;
wire w_0481_;
wire w_0482_;
wire w_0483_;
wire w_0484_;
wire w_0485_;
wire w_0486_;
wire w_0487_;
wire w_0488_;
wire w_0489_;
wire w_0490_;
wire w_0491_;
wire w_0492_;
wire w_0493_;
wire w_0494_;
wire w_0495_;
wire w_0496_;
wire w_0497_;
wire w_0498_;
wire w_0499_;
wire w_0500_;
wire w_0501_;
wire w_0502_;
wire w_0503_;
wire w_0504_;
wire w_0505_;
wire w_0506_;
wire w_0507_;
wire w_0508_;
wire w_0509_;
wire w_0510_;
wire w_0511_;
wire w_0512_;
wire w_0513_;
wire w_0514_;
wire w_0515_;
wire w_0516_;
wire w_0517_;
wire w_0518_;
wire w_0519_;
wire w_0520_;
wire w_0521_;
wire w_0522_;
wire w_0523_;
wire w_0524_;
wire w_0525_;
wire w_0526_;
wire w_0527_;
wire w_0528_;
wire w_0529_;
wire w_0530_;
wire w_0531_;
wire w_0532_;
wire w_0533_;
wire w_0534_;
wire w_0535_;
wire w_0536_;
wire w_0537_;
wire w_0538_;
wire w_0539_;
wire w_0540_;
wire w_0541_;
wire w_0542_;
wire w_0543_;
wire w_0544_;
wire w_0545_;
wire w_0546_;
wire w_0547_;
wire w_0548_;
wire w_0549_;
wire w_0550_;
wire w_0551_;
wire w_0552_;
wire w_0553_;
wire w_0554_;
wire w_0555_;
wire w_0556_;
wire w_0557_;
wire w_0558_;
wire w_0559_;
wire w_0560_;
wire w_0561_;
wire w_0562_;
wire w_0563_;
wire w_0564_;
wire w_0565_;
wire w_0566_;
wire w_0567_;
wire w_0568_;
wire w_0569_;
wire w_0570_;
wire w_0571_;
wire w_0572_;
wire w_0573_;
wire w_0574_;
wire w_0575_;
wire w_0576_;
wire w_0577_;
wire w_0578_;
wire w_0579_;
wire w_0580_;
wire w_0581_;
wire w_0582_;
wire w_0583_;
wire w_0584_;
wire w_0585_;
wire w_0586_;
wire w_0587_;
wire w_0588_;
wire w_0589_;
wire w_0590_;
wire w_0591_;
wire w_0592_;
wire w_0593_;
wire w_0594_;
wire w_0595_;
wire w_0596_;
wire w_0597_;
wire w_0598_;
wire w_0599_;
wire w_0600_;
wire w_0601_;
wire w_0602_;
wire w_0603_;
wire w_0604_;
wire w_0605_;
wire w_0606_;
wire w_0607_;
wire w_0608_;
wire w_0609_;
wire w_0610_;
wire w_0611_;
wire w_0612_;
wire w_0613_;
wire w_0614_;
wire w_0615_;
wire w_0616_;
wire w_0617_;
wire w_0618_;
wire w_0619_;
wire w_0620_;
wire w_0621_;
wire w_0622_;
wire w_0623_;
wire w_0624_;
wire w_0625_;
wire w_0626_;
wire w_0627_;
wire w_0628_;
wire w_0629_;
wire w_0630_;
wire w_0631_;
wire w_0632_;
wire w_0633_;
wire w_0634_;
wire w_0635_;
wire w_0636_;
wire w_0637_;
wire w_0638_;
wire w_0639_;
wire w_0640_;
wire w_0641_;
wire w_0642_;
wire w_0643_;
wire w_0644_;
wire w_0645_;
wire w_0646_;
wire w_0647_;
wire w_0648_;
wire w_0649_;
wire w_0650_;
wire w_0651_;
wire w_0652_;
wire w_0653_;
wire w_0654_;
wire w_0655_;
wire w_0656_;
wire w_0657_;
wire w_0658_;
wire w_0659_;
wire w_0660_;
wire w_0661_;
wire w_0662_;
wire w_0663_;
wire w_0664_;
wire w_0665_;
wire w_0666_;
wire w_0667_;
wire w_0668_;
wire w_0669_;
wire w_0670_;
wire w_0671_;
wire w_0672_;
wire w_0673_;
wire w_0674_;
wire w_0675_;
wire w_0676_;
wire w_0677_;
wire w_0678_;
wire w_0679_;
wire w_0680_;
wire w_0681_;
wire w_0682_;
wire w_0683_;
wire w_0684_;
wire w_0685_;
wire w_0686_;
wire w_0687_;
wire w_0688_;
wire w_0689_;
wire w_0690_;
wire w_0691_;
wire w_0692_;
wire w_0693_;
wire w_0694_;
wire w_0695_;
wire w_0696_;
wire w_0697_;
wire w_0698_;
wire w_0699_;
wire w_0700_;
wire w_0701_;
wire w_0702_;
wire w_0703_;
wire w_0704_;
wire w_0705_;
wire w_0706_;
wire w_0707_;
wire w_0708_;
wire w_0709_;
wire w_0710_;
wire w_0711_;
wire w_0712_;
wire w_0713_;
wire w_0714_;
wire w_0715_;
wire w_0716_;
wire w_0717_;
wire w_0718_;
wire w_0719_;
wire w_0720_;
wire w_0721_;
wire w_0722_;
wire w_0723_;
wire w_0724_;
wire w_0725_;
wire w_0726_;
wire w_0727_;
wire w_0728_;
wire w_0729_;
wire w_0730_;
wire w_0731_;
wire w_0732_;
wire w_0733_;
wire w_0734_;
wire w_0735_;
wire w_0736_;
wire w_0737_;
wire w_0738_;
wire w_0739_;
wire w_0740_;
wire w_0741_;
wire w_0742_;
wire w_0743_;
wire w_0744_;
wire w_0745_;
wire w_0746_;
wire w_0747_;
wire w_0748_;
wire w_0749_;
wire w_0750_;
wire w_0751_;
wire w_0752_;
wire w_0753_;
wire w_0754_;
wire w_0755_;
wire w_0756_;
wire w_0757_;
wire w_0758_;
wire w_0759_;
wire w_0760_;
wire w_0761_;
wire w_0762_;
wire w_0763_;
wire w_0764_;
wire w_0765_;
wire w_0766_;
wire w_0767_;
wire w_0768_;
wire w_0769_;
wire w_0770_;
wire w_0771_;
wire w_0772_;
wire w_0773_;
wire w_0774_;
wire w_0775_;
wire w_0776_;
wire w_0777_;
wire w_0778_;
wire w_0779_;
wire w_0780_;
wire w_0781_;
wire w_0782_;
wire w_0783_;
wire w_0784_;
wire w_0785_;
wire w_0786_;
wire w_0787_;
wire w_0788_;
wire w_0789_;
wire w_0790_;
wire w_0791_;
wire w_0792_;
wire w_0793_;
wire w_0794_;
wire w_0795_;
wire w_0796_;
wire w_0797_;
wire w_0798_;
wire w_0799_;
wire w_0800_;
wire w_0801_;
wire w_0802_;
wire w_0803_;
wire w_0804_;
wire w_0805_;
wire w_0806_;
wire w_0807_;
wire w_0808_;
wire w_0809_;
wire w_0810_;
wire w_0811_;
wire w_0812_;
wire w_0813_;
wire w_0814_;
wire w_0815_;
wire w_0816_;
wire w_0817_;
wire w_0818_;
wire w_0819_;
wire w_0820_;
wire w_0821_;
wire w_0822_;
wire w_0823_;
wire w_0824_;
wire w_0825_;
wire w_0826_;
wire w_0827_;
wire w_0828_;
wire w_0829_;
wire w_0830_;
wire w_0831_;
wire w_0832_;
wire w_0833_;
wire w_0834_;
wire w_0835_;
wire w_0836_;
wire w_0837_;
wire w_0838_;
wire w_0839_;
wire w_0840_;
wire w_0841_;
wire w_0842_;
wire w_0843_;
wire w_0844_;
wire w_0845_;
wire w_0846_;
wire w_0847_;
wire w_0848_;
wire w_0849_;
wire w_0850_;
wire w_0851_;
wire w_0852_;
wire w_0853_;
wire w_0854_;
wire w_0855_;
wire w_0856_;
wire w_0857_;
wire w_0858_;
wire w_0859_;
wire w_0860_;
wire w_0861_;
wire w_0862_;
wire w_0863_;
wire w_0864_;
wire w_0865_;
wire w_0866_;
wire w_0867_;
wire w_0868_;
wire w_0869_;
wire w_0870_;
wire w_0871_;
wire w_0872_;
wire w_0873_;
wire w_0874_;
wire w_0875_;
wire w_0876_;
wire w_0877_;
wire w_0878_;
wire w_0879_;
wire w_0880_;
wire w_0881_;
wire w_0882_;
wire w_0883_;
wire w_0884_;
wire w_0885_;
wire w_0886_;
wire w_0887_;
wire w_0888_;
wire w_0889_;
wire w_0890_;
wire w_0891_;
wire w_0892_;
wire w_0893_;
wire w_0894_;
wire w_0895_;
wire w_0896_;
wire w_0897_;
wire w_0898_;
wire w_0899_;
wire w_0900_;
wire w_0901_;
wire w_0902_;
wire w_0903_;
wire w_0904_;
wire w_0905_;
wire w_0906_;
wire w_0907_;
wire w_0908_;
wire w_0909_;
wire w_0910_;
wire w_0911_;
wire w_0912_;
wire w_0913_;
wire w_0914_;
wire w_0915_;
wire w_0916_;
wire w_0917_;
wire w_0918_;
wire w_0919_;
wire w_0920_;
wire w_0921_;
wire w_0922_;
wire w_0923_;
wire w_0924_;
wire w_0925_;
wire w_0926_;
wire w_0927_;
wire w_0928_;
wire w_0929_;
wire w_0930_;
wire w_0931_;
wire w_0932_;
wire w_0933_;
wire w_0934_;
wire w_0935_;
wire w_0936_;
wire w_0937_;
wire w_0938_;
wire w_0939_;
wire w_0940_;
wire w_0941_;
wire w_0942_;
wire w_0943_;
wire w_0944_;
wire w_0945_;
wire w_0946_;
wire w_0947_;
wire w_0948_;
wire w_0949_;
wire w_0950_;
wire w_0951_;
wire w_0952_;
wire w_0953_;
wire w_0954_;
wire w_0955_;
wire w_0956_;
wire w_0957_;
wire w_0958_;
wire w_0959_;
wire w_0960_;
wire w_0961_;
wire w_0962_;
wire w_0963_;
wire w_0964_;
wire w_0965_;
wire w_0966_;
wire w_0967_;
wire w_0968_;
wire w_0969_;
wire w_0970_;
wire w_0971_;
wire w_0972_;
wire w_0973_;
wire w_0974_;
wire w_0975_;
wire w_0976_;
wire w_0977_;
wire w_0978_;
wire w_0979_;
wire w_0980_;
wire w_0981_;
wire w_0982_;
wire w_0983_;
wire w_0984_;
wire w_0985_;
wire w_0986_;
wire w_0987_;
wire w_0988_;
wire w_0989_;
wire w_0990_;
wire w_0991_;
wire w_0992_;
wire w_0993_;
wire w_0994_;
wire w_0995_;
wire w_0996_;
wire w_0997_;
wire w_0998_;
wire w_0999_;
wire w_1000_;
wire w_1001_;
wire w_1002_;
wire w_1003_;
wire w_1004_;
wire w_1005_;
wire w_1006_;
wire w_1007_;
wire w_1008_;
wire w_1009_;
wire w_1010_;
wire w_1011_;
wire w_1012_;
wire w_1013_;
wire w_1014_;
wire w_1015_;
wire w_1016_;
wire w_1017_;
wire w_1018_;
wire w_1019_;
wire w_1020_;
wire w_1021_;
wire w_1022_;
wire w_1023_;
wire w_1024_;
wire w_1025_;
wire w_1026_;
wire w_1027_;
wire w_1028_;
wire w_1029_;
wire w_1030_;
wire w_1031_;
wire w_1032_;
wire w_1033_;
wire w_1034_;
wire w_1035_;
wire w_1036_;
wire w_1037_;
wire w_1038_;
wire w_1039_;
wire w_1040_;
wire w_1041_;
wire w_1042_;
wire w_1043_;
wire w_1044_;
wire w_1045_;
wire w_1046_;
wire w_1047_;
wire w_1048_;
wire w_1049_;
wire w_1050_;
wire w_1051_;
wire w_1052_;
wire w_1053_;
wire w_1054_;
wire w_1055_;
wire w_1056_;
wire w_1057_;
wire w_1058_;
wire w_1059_;
wire w_1060_;
wire w_1061_;
wire w_1062_;
wire w_1063_;
wire w_1064_;
wire w_1065_;
wire w_1066_;
wire w_1067_;
wire w_1068_;
wire w_1069_;
wire w_1070_;
wire w_1071_;
wire w_1072_;
wire w_1073_;
wire w_1074_;
wire w_1075_;
wire w_1076_;
wire w_1077_;
wire w_1078_;
wire w_1079_;
wire w_1080_;
wire w_1081_;
wire w_1082_;
wire w_1083_;
wire w_1084_;
wire w_1085_;
wire w_1086_;
wire w_1087_;
wire w_1088_;
wire w_1089_;
wire w_1090_;
wire w_1091_;
wire w_1092_;
wire w_1093_;
wire w_1094_;
wire w_1095_;
wire w_1096_;
wire w_1097_;
wire w_1098_;
wire w_1099_;
wire w_1100_;
wire w_1101_;
wire w_1102_;
wire w_1103_;
wire w_1104_;
wire w_1105_;
wire w_1106_;
wire w_1107_;
wire w_1108_;
wire w_1109_;
wire w_1110_;
wire w_1111_;
wire w_1112_;
wire w_1113_;
wire w_1114_;
wire w_1115_;
wire w_1116_;
wire w_1117_;
wire w_1118_;
wire w_1119_;
wire w_1120_;
wire w_1121_;
wire w_1122_;
wire w_1123_;
wire w_1124_;
wire w_1125_;
wire w_1126_;
wire w_1127_;
wire w_1128_;
wire w_1129_;
wire w_1130_;
wire w_1131_;
wire w_1132_;
wire w_1133_;
wire w_1134_;
wire w_1135_;
wire w_1136_;
wire w_1137_;
wire w_1138_;
wire w_1139_;
wire w_1140_;
wire w_1141_;
wire w_1142_;
wire w_1143_;
wire w_1144_;
wire w_1145_;
wire w_1146_;
wire w_1147_;
wire w_1148_;
wire w_1149_;
wire w_1150_;
wire w_1151_;
wire w_1152_;
wire w_1153_;
wire w_1154_;
wire w_1155_;
wire w_1156_;
wire w_1157_;
wire w_1158_;
wire w_1159_;
wire w_1160_;
wire w_1161_;
wire w_1162_;
wire w_1163_;
wire w_1164_;
wire w_1165_;
wire w_1166_;
wire w_1167_;
wire w_1168_;
wire w_1169_;
wire w_1170_;
wire w_1171_;
wire w_1172_;
wire w_1173_;
wire w_1174_;
wire w_1175_;
wire w_1176_;
wire w_1177_;
wire w_1178_;
wire w_1179_;
wire w_1180_;
wire w_1181_;
wire w_1182_;
wire w_1183_;
wire w_1184_;
wire w_1185_;
wire w_1186_;
wire w_1187_;
wire w_1188_;
wire w_1189_;
wire w_1190_;
wire w_1191_;
wire w_1192_;
wire w_1193_;
wire w_1194_;
wire w_1195_;
wire w_1196_;
wire w_1197_;
wire w_1198_;
wire w_1199_;
wire w_1200_;
wire w_1201_;
wire w_1202_;
wire w_1203_;
wire w_1204_;
wire w_1205_;
wire w_1206_;
wire w_1207_;
wire w_1208_;
wire w_1209_;
wire w_1210_;
wire w_1211_;
wire w_1212_;
wire w_1213_;
wire w_1214_;
wire w_1215_;
wire w_1216_;
wire w_1217_;
wire w_1218_;
wire w_1219_;
wire w_1220_;
wire w_1221_;
wire w_1222_;
wire w_1223_;
wire w_1224_;
wire w_1225_;
wire w_1226_;
wire w_1227_;
wire w_1228_;
wire w_1229_;
wire w_1230_;
wire w_1231_;
wire w_1232_;
wire w_1233_;
wire w_1234_;
wire w_1235_;
wire w_1236_;
wire w_1237_;
wire w_1238_;
wire w_1239_;
wire w_1240_;
wire w_1241_;
wire w_1242_;
wire w_1243_;
wire w_1244_;
wire w_1245_;
wire w_1246_;
wire w_1247_;
wire w_1248_;
wire w_1249_;
wire w_1250_;
wire w_1251_;
wire w_1252_;
wire w_1253_;
wire w_1254_;
wire w_1255_;
wire w_1256_;
wire w_1257_;
wire w_1258_;
wire w_1259_;
wire w_1260_;
wire w_1261_;
wire w_1262_;
wire w_1263_;
wire w_1264_;
wire w_1265_;
wire w_1266_;
wire w_1267_;
wire w_1268_;
wire w_1269_;
wire w_1270_;
wire w_1271_;
wire w_1272_;
wire w_1273_;
wire w_1274_;
wire w_1275_;
wire w_1276_;
wire w_1277_;
wire w_1278_;
wire w_1279_;
wire w_1280_;
wire w_1281_;
wire w_1282_;
wire w_1283_;
wire w_1284_;
wire w_1285_;
wire w_1286_;
wire w_1287_;
wire w_1288_;
wire w_1289_;
wire w_1290_;
wire w_1291_;
wire w_1292_;
wire w_1293_;
wire w_1294_;
wire w_1295_;
wire w_1296_;
wire w_1297_;
wire w_1298_;
wire w_1299_;
wire w_1300_;
wire w_1301_;
wire w_1302_;
wire w_1303_;
wire w_1304_;
wire w_1305_;
wire w_1306_;
wire w_1307_;
wire w_1308_;
wire w_1309_;
wire w_1310_;
wire w_1311_;
wire w_1312_;
wire w_1313_;
wire w_1314_;
wire w_1315_;
wire w_1316_;
wire w_1317_;
wire w_1318_;
wire w_1319_;
wire w_1320_;
wire w_1321_;
wire w_1322_;
wire w_1323_;
wire w_1324_;
wire w_1325_;
wire w_1326_;
wire w_1327_;
wire w_1328_;
wire w_1329_;
wire w_1330_;
wire w_1331_;
wire w_1332_;
wire w_1333_;
wire w_1334_;
wire w_1335_;
wire w_1336_;
wire w_1337_;
wire w_1338_;
wire w_1339_;
wire w_1340_;
wire w_1341_;
wire w_1342_;
wire w_1343_;
wire w_1344_;
wire w_1345_;
wire w_1346_;
wire w_1347_;
wire w_1348_;
wire w_1349_;
wire w_1350_;
wire w_1351_;
wire w_1352_;
wire w_1353_;
wire w_1354_;
wire w_1355_;
wire w_1356_;
wire w_1357_;
wire w_1358_;
wire w_1359_;
wire w_1360_;
wire w_1361_;
wire w_1362_;
wire w_1363_;
wire w_1364_;
wire w_1365_;
wire w_1366_;
wire w_1367_;
wire w_1368_;
wire w_1369_;
wire w_1370_;
wire w_1371_;
wire w_1372_;
wire w_1373_;
wire w_1374_;
wire w_1375_;
wire w_1376_;
wire w_1377_;
wire w_1378_;
wire w_1379_;
wire w_1380_;
wire w_1381_;
wire w_1382_;
wire w_1383_;
wire w_1384_;
wire w_1385_;
wire w_1386_;
wire w_1387_;
wire w_1388_;
wire w_1389_;
wire w_1390_;
wire w_1391_;
wire w_1392_;
wire w_1393_;
wire w_1394_;
wire w_1395_;
wire w_1396_;
wire w_1397_;
wire w_1398_;
wire w_1399_;
wire w_1400_;
wire w_1401_;
wire w_1402_;
wire w_1403_;
wire w_1404_;
wire w_1405_;
wire w_1406_;
wire w_1407_;
wire w_1408_;
wire w_1409_;
wire w_1410_;
wire w_1411_;
wire w_1412_;
wire w_1413_;
wire w_1414_;
wire w_1415_;
wire w_1416_;
wire w_1417_;
wire w_1418_;
wire w_1419_;
wire w_1420_;
wire w_1421_;
wire w_1422_;
wire w_1423_;
wire w_1424_;
wire w_1425_;
wire w_1426_;
wire w_1427_;
wire w_1428_;
wire w_1429_;
wire w_1430_;
wire w_1431_;
wire w_1432_;
wire w_1433_;
wire w_1434_;
wire w_1435_;
wire w_1436_;
wire w_1437_;
wire w_1438_;
wire w_1439_;
wire w_1440_;
wire w_1441_;
wire w_1442_;
wire w_1443_;
wire w_1444_;
wire w_1445_;
wire w_1446_;
wire w_1447_;
wire w_1448_;
wire w_1449_;
wire w_1450_;
wire w_1451_;
wire w_1452_;
wire w_1453_;
wire w_1454_;
wire w_1455_;
wire w_1456_;
wire w_1457_;
wire w_1458_;
wire w_1459_;
wire w_1460_;
wire w_1461_;
wire w_1462_;
wire w_1463_;
wire w_1464_;
wire w_1465_;
wire w_1466_;
wire w_1467_;
wire w_1468_;
wire w_1469_;
wire w_1470_;
wire w_1471_;
wire w_1472_;
wire w_1473_;
wire w_1474_;
wire w_1475_;
wire w_1476_;
wire w_1477_;
wire w_1478_;
wire w_1479_;
wire w_1480_;
wire w_1481_;
wire w_1482_;
wire w_1483_;
wire w_1484_;
wire w_1485_;
wire w_1486_;
wire w_1487_;
wire w_1488_;
wire w_1489_;
wire w_1490_;
wire w_1491_;
wire w_1492_;
wire w_1493_;
wire w_1494_;
wire w_1495_;
wire w_1496_;
wire w_1497_;
wire w_1498_;
wire w_1499_;
wire w_1500_;
wire w_1501_;
wire w_1502_;
wire w_1503_;
wire w_1504_;
wire w_1505_;
wire w_1506_;
wire w_1507_;
wire w_1508_;
wire w_1509_;
wire w_1510_;
wire w_1511_;
wire w_1512_;
wire w_1513_;
wire w_1514_;
wire w_1515_;
wire w_1516_;
wire w_1517_;
wire w_1518_;
wire w_1519_;
wire w_1520_;
wire w_1521_;
wire w_1522_;
wire w_1523_;
wire w_1524_;
wire w_1525_;
wire w_1526_;
wire w_1527_;
wire w_1528_;
wire w_1529_;
wire w_1530_;
wire w_1531_;
wire w_1532_;
wire w_1533_;
wire w_1534_;
wire w_1535_;
wire w_1536_;
wire w_1537_;
wire w_1538_;
wire w_1539_;
wire w_1540_;
wire w_1541_;
wire w_1542_;
wire w_1543_;
wire w_1544_;
wire w_1545_;
wire w_1546_;
wire w_1547_;
wire w_1548_;
wire w_1549_;
wire w_1550_;
wire w_1551_;
wire w_1552_;
wire w_1553_;
wire w_1554_;
wire w_1555_;
wire w_1556_;
wire w_1557_;
wire w_1558_;
wire w_1559_;
wire w_1560_;
wire w_1561_;
wire w_1562_;
wire w_1563_;
wire w_1564_;
wire w_1565_;
wire w_1566_;
wire w_1567_;
wire w_1568_;
wire w_1569_;
wire w_1570_;
wire w_1571_;
wire w_1572_;
wire w_1573_;
wire w_1574_;
wire w_1575_;
wire w_1576_;
wire w_1577_;
wire w_1578_;
wire w_1579_;
wire w_1580_;
wire w_1581_;
wire w_1582_;
wire w_1583_;
wire w_1584_;
wire w_1585_;
wire w_1586_;
wire w_1587_;
wire w_1588_;
wire w_1589_;
wire w_1590_;
wire w_1591_;
wire w_1592_;
wire w_1593_;
wire w_1594_;
wire w_1595_;
wire w_1596_;
wire w_1597_;
wire w_1598_;
wire w_1599_;
wire w_1600_;
wire w_1601_;
wire w_1602_;
wire w_1603_;
wire w_1604_;
wire w_1605_;
wire w_1606_;
wire w_1607_;
wire w_1608_;
wire w_1609_;
wire w_1610_;
wire w_1611_;
wire w_1612_;
wire w_1613_;
wire w_1614_;
wire w_1615_;
wire w_1616_;
wire w_1617_;
wire w_1618_;
wire w_1619_;
wire w_1620_;
wire w_1621_;
wire w_1622_;
wire w_1623_;
wire w_1624_;
wire w_1625_;
wire w_1626_;
wire w_1627_;
wire w_1628_;
wire w_1629_;
wire w_1630_;
wire w_1631_;
wire w_1632_;
wire w_1633_;
wire w_1634_;
wire w_1635_;
wire w_1636_;
wire w_1637_;
wire w_1638_;
wire w_1639_;
wire w_1640_;
wire w_1641_;
wire w_1642_;
wire w_1643_;
wire w_1644_;
wire w_1645_;
wire w_1646_;
wire w_1647_;
wire w_1648_;
wire w_1649_;
wire w_1650_;
wire w_1651_;
wire w_1652_;
wire w_1653_;
wire w_1654_;
wire w_1655_;
wire w_1656_;
wire w_1657_;
wire w_1658_;
wire w_1659_;
wire w_1660_;
wire w_1661_;
wire w_1662_;
wire w_1663_;
wire w_1664_;
wire w_1665_;
wire w_1666_;
wire w_1667_;
wire w_1668_;
wire w_1669_;
wire w_1670_;
wire w_1671_;
wire w_1672_;
wire w_1673_;
wire w_1674_;
wire w_1675_;
wire w_1676_;
wire w_1677_;
wire w_1678_;
wire w_1679_;
wire w_1680_;
wire w_1681_;
wire w_1682_;
wire w_1683_;
wire w_1684_;
wire w_1685_;
wire w_1686_;
wire w_1687_;
wire w_1688_;
wire w_1689_;
wire w_1690_;
wire w_1691_;
wire w_1692_;
wire w_1693_;
wire w_1694_;
wire w_1695_;
wire w_1696_;
wire w_1697_;
wire w_1698_;
wire w_1699_;
wire w_1700_;
wire w_1701_;
wire w_1702_;
wire w_1703_;
wire w_1704_;
wire w_1705_;
wire w_1706_;
wire w_1707_;
wire w_1708_;
wire w_1709_;
wire w_1710_;
wire w_1711_;
wire w_1712_;
wire w_1713_;
wire w_1714_;
wire w_1715_;
wire w_1716_;
wire w_1717_;
wire w_1718_;
wire w_1719_;
wire w_1720_;
wire w_1721_;
wire w_1722_;
wire w_1723_;
wire w_1724_;
wire w_1725_;
wire w_1726_;
wire w_1727_;
wire w_1728_;
wire w_1729_;
wire w_1730_;
wire w_1731_;
wire w_1732_;
wire w_1733_;
wire w_1734_;
wire w_1735_;
wire w_1736_;
wire w_1737_;
wire w_1738_;
wire w_1739_;
wire w_1740_;
wire w_1741_;
wire w_1742_;
wire w_1743_;
wire w_1744_;
wire w_1745_;
wire w_1746_;
wire w_1747_;
wire w_1748_;
wire w_1749_;
wire w_1750_;
wire w_1751_;
wire w_1752_;
wire w_1753_;
wire w_1754_;
wire w_1755_;
wire w_1756_;
wire w_1757_;
wire w_1758_;
wire w_1759_;
wire w_1760_;
wire w_1761_;
wire w_1762_;
wire w_1763_;
wire w_1764_;
wire w_1765_;
wire w_1766_;
wire w_1767_;
wire w_1768_;
wire w_1769_;
wire w_1770_;
wire w_1771_;
wire w_1772_;
wire w_1773_;
wire w_1774_;
wire w_1775_;
wire w_1776_;
wire w_1777_;
wire w_1778_;
wire w_1779_;
wire w_1780_;
wire w_1781_;
wire w_1782_;
wire w_1783_;
wire w_1784_;
wire w_1785_;
wire w_1786_;
wire w_1787_;
wire w_1788_;
wire w_1789_;
wire w_1790_;
wire w_1791_;
wire w_1792_;
wire w_1793_;
wire w_1794_;
wire w_1795_;
wire w_1796_;
wire w_1797_;
wire w_1798_;
wire w_1799_;
wire w_1800_;
wire w_1801_;
wire w_1802_;
wire w_1803_;
wire w_1804_;
wire w_1805_;
wire w_1806_;
wire w_1807_;
wire w_1808_;
wire w_1809_;
wire w_1810_;
wire w_1811_;
wire w_1812_;
wire w_1813_;
wire w_1814_;
wire w_1815_;
wire w_1816_;
wire w_1817_;
wire w_1818_;
wire w_1819_;
wire w_1820_;
wire w_1821_;
wire w_1822_;
wire w_1823_;
wire w_1824_;
wire w_1825_;
wire w_1826_;
wire w_1827_;
wire w_1828_;
wire w_1829_;
wire w_1830_;
wire w_1831_;
wire w_1832_;
wire w_1833_;
wire w_1834_;
wire w_1835_;
wire w_1836_;
wire w_1837_;
wire w_1838_;
wire w_1839_;
wire w_1840_;
wire w_1841_;
wire w_1842_;
wire w_1843_;
wire w_1844_;
wire w_1845_;
wire w_1846_;
wire w_1847_;
wire w_1848_;
wire w_1849_;
wire w_1850_;
wire w_1851_;
wire w_1852_;
wire w_1853_;
wire w_1854_;
wire w_1855_;
wire w_1856_;
wire w_1857_;
wire w_1858_;
wire w_1859_;
wire w_1860_;
wire w_1861_;
wire w_1862_;
wire w_1863_;
wire w_1864_;
wire w_1865_;
wire w_1866_;
wire w_1867_;
wire w_1868_;
wire w_1869_;
wire w_1870_;
wire w_1871_;
wire w_1872_;
wire w_1873_;
wire w_1874_;
wire w_1875_;
wire w_1876_;
wire w_1877_;
wire w_1878_;
wire w_1879_;
wire w_1880_;
wire w_1881_;
wire w_1882_;
wire w_1883_;
wire w_1884_;
wire w_1885_;
wire w_1886_;
wire w_1887_;
wire w_1888_;
wire w_1889_;
wire w_1890_;
wire w_1891_;
wire w_1892_;
wire w_1893_;
wire w_1894_;
wire w_1895_;
wire w_1896_;
wire w_1897_;
wire w_1898_;
wire w_1899_;
wire w_1900_;
wire w_1901_;
wire w_1902_;
wire w_1903_;
wire w_1904_;
wire w_1905_;
wire w_1906_;
wire w_1907_;
wire w_1908_;
wire w_1909_;
wire w_1910_;
wire w_1911_;
wire w_1912_;
wire w_1913_;
wire w_1914_;
wire w_1915_;
wire w_1916_;
wire w_1917_;
wire w_1918_;
wire w_1919_;
wire w_1920_;
wire w_1921_;
wire w_1922_;
wire w_1923_;
wire w_1924_;
wire w_1925_;
wire w_1926_;
wire w_1927_;
wire w_1928_;
wire w_1929_;
wire w_1930_;
wire w_1931_;
wire w_1932_;
wire w_1933_;
wire w_1934_;
wire w_1935_;
wire w_1936_;
wire w_1937_;
wire w_1938_;
wire w_1939_;
wire w_1940_;
wire w_1941_;
wire w_1942_;
wire w_1943_;
wire w_1944_;
wire w_1945_;
wire w_1946_;
wire w_1947_;
wire w_1948_;
wire w_1949_;
wire w_1950_;
wire w_1951_;
wire w_1952_;
wire w_1953_;
wire w_1954_;
wire w_1955_;
wire w_1956_;
wire w_1957_;
wire w_1958_;
wire w_1959_;
wire w_1960_;
wire w_1961_;
wire w_1962_;
wire w_1963_;
wire w_1964_;
wire w_1965_;
wire w_1966_;
wire w_1967_;
wire w_1968_;
wire w_1969_;
wire w_1970_;
wire w_1971_;
wire w_1972_;
wire w_1973_;
wire w_1974_;
wire w_1975_;
wire w_1976_;
wire w_1977_;
wire w_1978_;
wire w_1979_;
wire w_1980_;
wire w_1981_;
wire w_1982_;
wire w_1983_;
wire w_1984_;
wire w_1985_;
wire w_1986_;
wire w_1987_;
wire w_1988_;
wire w_1989_;
wire w_1990_;
wire w_1991_;
wire w_1992_;
wire w_1993_;
wire w_1994_;
wire w_1995_;
wire w_1996_;
wire w_1997_;
wire w_1998_;
wire w_1999_;
wire w_2000_;
wire w_2001_;
wire w_2002_;
wire w_2003_;
wire w_2004_;
wire w_2005_;
wire w_2006_;
wire w_2007_;
wire w_2008_;
wire w_2009_;
wire w_2010_;
wire w_2011_;
wire w_2012_;
wire w_2013_;
wire w_2014_;
wire w_2015_;
wire w_2016_;
wire w_2017_;
wire w_2018_;
wire w_2019_;
wire w_2020_;
wire w_2021_;
wire w_2022_;
wire w_2023_;
wire w_2024_;
wire w_2025_;
wire w_2026_;
wire w_2027_;
wire w_2028_;
wire w_2029_;
wire w_2030_;
wire w_2031_;
wire w_2032_;
wire w_2033_;
wire w_2034_;
wire w_2035_;
wire w_2036_;
wire w_2037_;
wire w_2038_;
wire w_2039_;
wire w_2040_;
wire w_2041_;
wire w_2042_;
wire w_2043_;
wire w_2044_;
wire w_2045_;
wire w_2046_;
wire w_2047_;
wire w_2048_;
wire w_2049_;
wire w_2050_;
wire w_2051_;
wire w_2052_;
wire w_2053_;
wire w_2054_;
wire w_2055_;
wire w_2056_;
wire w_2057_;
wire w_2058_;
wire w_2059_;
wire w_2060_;
wire w_2061_;
wire w_2062_;
wire w_2063_;
wire w_2064_;
wire w_2065_;
wire w_2066_;
wire w_2067_;
wire w_2068_;
wire w_2069_;
wire w_2070_;
wire w_2071_;
wire w_2072_;
wire w_2073_;
wire w_2074_;
wire w_2075_;
wire w_2076_;
wire w_2077_;
wire w_2078_;
wire w_2079_;
wire w_2080_;
wire w_2081_;
wire w_2082_;
wire w_2083_;
wire w_2084_;
wire w_2085_;
wire w_2086_;
wire w_2087_;
wire w_2088_;
wire w_2089_;
wire w_2090_;
wire w_2091_;
wire w_2092_;
wire w_2093_;
wire w_2094_;
wire w_2095_;
wire w_2096_;
wire w_2097_;
wire w_2098_;
wire w_2099_;
xor (w_1438_, w_1435_, w_0528_);
nand (w_0036_, new_in5[3], new_in2[3]);
and (w_1455_, new_in6[1], new_in10[5]);
and (w_1302_, w_1067_, w_1975_);
nand (w_2094_, w_1103_, w_0193_);
nand (new_out8[3], w_1307_, w_1335_);
xor (w_0904_, new_in5[1], new_in2[0]);
xor (w_0603_, w_0958_, w_0096_);
or (w_1062_, w_1896_, w_0807_);
nand (w_1570_, w_1704_, w_0759_);
xor (w_0935_, w_1337_, w_0298_);
nand (w_1090_, w_1708_, w_0073_);
nand (w_1019_, w_0493_, w_0809_);
xor (w_2091_, w_1317_, w_1610_);
xor (w_1001_, new_in11[0], new_in7[0]);
and (new_out11[2], w_0200_, w_0427_);
and (w_1088_, w_1585_, w_0794_);
and (w_1728_, new_in1[2], new_in3[1]);
xor (w_1262_, w_0410_, w_1659_);
nand (w_1205_, w_0565_, w_2006_);
nand (w_0397_, w_1398_, w_0663_);
nand (w_0097_, new_in2[6], new_in6[4]);
and (w_0205_, new_in5[1], new_in2[0]);
nand (w_0206_, w_0045_, w_1330_);
nand (w_0676_, w_1650_, w_0011_);
nand (w_2047_, new_in8[1], new_in3[1]);
xor (w_0545_, new_in6[4], new_in4[4]);
nand (w_1133_, w_0802_, w_1239_);
and (w_2096_, w_1931_, w_1233_);
xor (w_1305_, new_in10[2], w_1416_);
and (w_0788_, new_in10[3], new_in4[6]);
nand (w_1606_, w_0200_, w_0693_);
xor (w_1998_, w_1952_, w_2026_);
nand (w_2025_, w_0638_, w_0089_);
not (w_1817_, w_0730_);
and (w_1181_, new_in11[0], new_in7[0]);
nand (w_0590_, w_1857_, w_1438_);
nand (w_1039_, w_1642_, w_2075_);
xor (w_0480_, w_1941_, w_0173_);
nand (w_2098_, w_1708_, w_0154_);
and (w_0031_, w_1244_, w_0341_);
nand (w_0091_, w_1679_, w_0247_);
and (w_0514_, w_0978_, w_1081_);
and (w_0309_, w_0217_, w_1184_);
xor (w_1634_, w_0479_, w_1792_);
xor (w_1555_, new_in4[8], new_in6[8]);
nand (w_0734_, w_1548_, w_1982_);
xor (w_1904_, w_0702_, w_0382_);
xor (w_1356_, w_1483_, w_1169_);
nand (w_1022_, new_in5[7], new_in3[4]);
nand (w_1971_, w_1985_, w_1655_);
xor (w_2097_, w_1533_, w_1214_);
nand (w_1292_, w_0217_, w_0328_);
xor (w_0813_, w_1734_, w_0988_);
nand (w_1778_, w_1857_, w_0362_);
and (w_1464_, new_in1[1], new_in3[3]);
xor (w_0773_, w_0377_, w_0042_);
nand (w_1824_, w_0318_, w_1622_);
xor (w_0141_, w_1513_, w_1953_);
nand (w_1100_, w_2028_, w_0907_);
xor (w_1320_, new_in5[0], new_in10[0]);
nand (w_1541_, w_1142_, w_0235_);
and (w_0954_, new_in1[1], new_in3[1]);
or (w_0202_, w_0189_, w_1842_);
nand (w_1535_, w_0041_, w_0024_);
nand (w_0538_, w_1181_, w_0846_);
and (w_1157_, new_in6[1], w_1999_);
xor (w_0876_, new_in2[3], w_0780_);
xor (w_1637_, new_in6[6], new_in2[1]);
xor (w_0696_, new_in8[3], new_in4[5]);
nand (w_1994_, w_1839_, w_0407_);
xor (w_1588_, new_in10[0], new_in3[1]);
and (w_0189_, new_in11[0], w_0785_);
xor (w_1544_, w_1847_, w_0688_);
xor (w_2065_, w_1823_, w_1827_);
nand (w_0409_, w_1568_, w_1179_);
xor (w_1922_, w_0503_, w_0162_);
xor (w_0464_, w_1041_, w_0612_);
xor (w_0304_, new_in2[6], new_in6[2]);
xor (w_1857_, w_1485_, w_0144_);
nand (w_1401_, w_1857_, w_0481_);
xor (w_1859_, w_0142_, w_1399_);
xor (w_0712_, new_in3[0], w_2077_);
nand (w_0316_, w_1031_, w_1489_);
and (w_1983_, new_in6[0], new_in10[5]);
or (w_0109_, w_1827_, w_0732_);
nand (w_1720_, w_1473_, w_1654_);
xor (w_0754_, new_in6[6], new_in7[1]);
and (w_1814_, w_0522_, w_1421_);
nand (w_0319_, new_in3[1], new_in2[2]);
xor (w_0659_, w_0864_, w_1346_);
and (w_0116_, new_in10[0], new_in7[0]);
xor (w_0847_, w_1888_, w_0195_);
nand (w_1840_, w_1183_, w_1553_);
xor (w_1595_, new_in8[2], w_1070_);
nand (new_out7[0], w_1970_, w_1865_);
xor (w_2014_, w_0367_, w_0941_);
nand (w_0708_, new_in6[6], new_in2[1]);
and (w_1160_, new_in10[2], new_in2[1]);
nand (w_0967_, w_0690_, w_1278_);
xor (w_0915_, w_1599_, w_0675_);
xor (w_0359_, w_0240_, w_0801_);
and (w_1473_, w_0958_, w_0096_);
xor (w_0850_, w_0378_, w_0550_);
nand (w_0908_, w_1453_, w_1955_);
or (w_0571_, w_0482_, w_1964_);
nand (w_1911_, w_1033_, w_1246_);
xor (w_1813_, w_1252_, w_0630_);
nand (w_0842_, w_1432_, w_0043_);
nand (w_0956_, w_0099_, w_0576_);
nand (w_1918_, w_0463_, w_1635_);
xor (w_1282_, new_in8[2], w_1227_);
or (w_1102_, w_0726_, w_1591_);
xor (w_1608_, w_1426_, new_in2[2]);
or (w_1023_, w_1708_, w_1369_);
xor (w_1920_, new_in10[2], w_0398_);
nand (w_1989_, w_1959_, w_1821_);
nand (w_1329_, w_0956_, w_0761_);
and (w_0416_, w_0425_, w_2018_);
xor (w_1761_, w_0295_, w_1457_);
and (w_0565_, new_in6[0], new_in2[2]);
and (w_1138_, w_2028_, w_0238_);
nand (w_0452_, w_1933_, w_0202_);
nand (w_1781_, w_0810_, w_0897_);
nand (w_1770_, w_0734_, w_1396_);
xor (w_1947_, w_1264_, w_1727_);
xor (w_1569_, new_in6[6], new_in5[2]);
xor (w_1797_, w_1142_, w_0235_);
xor (w_1846_, w_0325_, w_1728_);
xor (w_0761_, new_in8[2], new_in4[2]);
xor (w_0146_, new_in8[2], w_0291_);
xor (w_0724_, w_0700_, w_1886_);
and (w_1916_, new_in2[1], new_in5[3]);
nor (w_0674_, new_in8[2], new_in9[2]);
nand (w_0300_, w_0168_, w_1344_);
xor (w_0043_, w_1595_, w_1929_);
xor (w_1421_, w_1195_, w_0038_);
xor (w_2006_, new_in6[1], new_in2[3]);
xor (w_0253_, w_1053_, w_0850_);
nor (w_1155_, w_1406_, new_in1[2]);
xor (w_1733_, w_0030_, w_0696_);
nand (w_1311_, w_1038_, w_1468_);
and (w_1186_, new_in10[0], new_in4[0]);
nand (w_1389_, w_0168_, w_1077_);
nand (w_0102_, w_1548_, w_1141_);
xor (w_0107_, w_0828_, w_0118_);
nand (w_0308_, new_in6[2], new_in2[4]);
xor (w_0395_, w_1243_, w_1510_);
xor (w_0076_, new_in6[4], new_in5[3]);
nand (w_1388_, w_1715_, w_0392_);
and (w_1334_, w_0517_, w_0397_);
nand (w_1279_, w_0837_, w_0579_);
xor (w_2054_, w_1808_, w_2002_);
nand (w_1194_, w_0567_, w_0781_);
xor (w_0629_, w_0190_, w_1653_);
xor (w_1429_, w_1252_, new_in9[1]);
nand (new_out2, w_0699_, w_0859_);
xor (w_0444_, new_in6[5], new_in3[0]);
and (w_1783_, w_1632_, w_1493_);
and (w_0984_, new_in9[0], new_in8[1]);
xor (w_2003_, new_in3[1], w_1997_);
xor (w_0218_, w_1652_, w_1313_);
xor (w_1222_, new_in4[2], new_in5[6]);
and (w_0899_, w_1890_, w_0074_);
nand (w_1516_, w_0217_, w_1956_);
nand (w_1759_, w_0200_, w_1514_);
nand (w_1307_, w_0200_, w_1242_);
xor (w_0459_, w_1704_, w_0759_);
xor (w_0655_, w_0376_, w_1144_);
nand (new_out3[3], w_0647_, w_0604_);
nand (w_1109_, w_0959_, w_0776_);
xor (w_1384_, w_1107_, w_1156_);
or (w_1568_, w_0726_, w_1454_);
and (w_0642_, w_0810_, w_1340_);
xor (w_1332_, new_in8[3], new_in9[3]);
and (w_0408_, new_in2[3], new_in5[4]);
and (w_1518_, w_0983_, w_1275_);
nand (w_0871_, new_in3[2], new_in2[3]);
xor (w_1713_, w_1133_, w_1037_);
xor (w_1230_, w_1825_, w_0563_);
nand (w_0071_, w_0263_, w_1884_);
and (w_0227_, w_0266_, w_1414_);
xor (w_0376_, w_1669_, w_1064_);
and (w_0668_, w_2040_, w_0575_);
xor (w_0977_, w_0161_, w_1491_);
nand (w_0128_, w_0479_, w_0145_);
or (w_1621_, w_1705_, w_2065_);
nand (w_1527_, w_0488_, new_in6[2]);
xor (w_1373_, new_in5[2], new_in2[2]);
and (w_0487_, w_0133_, w_0534_);
nand (w_0586_, w_1752_, w_0181_);
nand (w_0684_, w_0276_, w_2061_);
xor (w_1950_, w_0230_, w_0119_);
nand (w_1269_, w_1833_, w_0433_);
xor (w_0435_, w_1976_, w_1336_);
nand (w_1868_, w_0747_, w_0892_);
xor (w_0342_, w_2005_, w_0009_);
nand (w_1263_, w_1708_, w_1717_);
xor (w_0127_, w_1890_, w_0074_);
xor (w_0414_, new_in6[3], w_0862_);
xor (w_1037_, new_in3[2], new_in2[2]);
xor (w_1313_, w_0870_, w_1464_);
xor (w_1547_, new_in10[3], w_0714_);
nand (w_0428_, w_0952_, w_1569_);
nand (w_1662_, w_1708_, w_1867_);
nand (w_1737_, w_1674_, w_0544_);
and (w_1104_, new_in8[3], new_in1[2]);
xor (w_0083_, w_0919_, w_0307_);
and (w_1636_, new_in8[1], new_in9[6]);
nand (w_0614_, w_0975_, w_0208_);
xor (w_0528_, w_0749_, w_0982_);
xor (w_0753_, new_in10[0], new_in6[0]);
nand (w_0736_, w_0726_, w_1950_);
nand (w_1985_, w_1834_, w_0039_);
xor (w_0010_, w_0368_, w_1905_);
and (w_1627_, w_1545_, w_0783_);
xor (w_1344_, w_1320_, w_0223_);
nand (new_out9[1], w_0869_, w_0406_);
nand (w_1562_, w_0151_, w_1481_);
nand (w_1832_, w_0846_, w_0058_);
xor (w_1066_, new_in6[1], w_1337_);
nand (w_0495_, w_0210_, w_0000_);
nand (w_0533_, w_1708_, w_0569_);
xor (w_0063_, w_1911_, w_0104_);
and (w_0118_, w_1295_, w_1226_);
and (w_1233_, new_in10[3], new_in3[1]);
and (w_0594_, w_1668_, w_0351_);
nand (w_1142_, w_2029_, w_1205_);
or (w_1200_, w_0726_, w_0923_);
nand (w_1533_, new_in10[3], new_in6[3]);
nand (w_0924_, w_1523_, w_0955_);
and (w_1005_, w_0760_, w_1304_);
nand (w_2040_, new_in6[1], w_1803_);
nand (w_0805_, w_1062_, w_1738_);
or (w_0470_, new_in5[1], w_1782_);
or (w_0451_, w_1825_, w_0563_);
nand (w_0577_, w_1708_, w_1562_);
and (w_0047_, w_1857_, w_0865_);
or (w_1521_, new_in5[0], w_0987_);
and (w_0216_, w_0560_, w_0131_);
nand (w_0510_, w_0372_, w_1091_);
nand (w_1703_, w_1360_, w_0265_);
nand (w_1440_, w_1931_, w_0726_);
and (w_0931_, w_0358_, w_1694_);
xor (w_1849_, w_1469_, w_0885_);
xor (w_0606_, w_2096_, w_0808_);
and (w_0556_, new_in8[3], new_in1[0]);
xor (w_1591_, new_in8[4], w_2046_);
xor (w_0130_, w_1034_, w_0805_);
nand (w_0479_, new_in9[0], new_in8[0]);
nand (w_0776_, w_0640_, w_1189_);
and (w_1546_, w_0913_, w_1858_);
nand (w_1322_, w_1857_, w_0074_);
xor (w_1220_, w_1816_, w_0607_);
nand (w_1903_, w_1597_, w_0856_);
or (w_1583_, w_0047_, w_0625_);
nand (w_1821_, w_1548_, w_0632_);
xor (w_0126_, w_1154_, w_1105_);
xor (w_1333_, w_0336_, w_1069_);
nand (w_2030_, w_1249_, w_0666_);
xor (w_1119_, new_in6[0], w_1337_);
or (w_0990_, w_0726_, w_2055_);
xor (w_2012_, w_0110_, w_0454_);
and (new_out1[0], w_0515_, w_0087_);
xor (w_1035_, w_1355_, w_0915_);
and (w_1910_, w_1104_, w_1466_);
nand (w_1902_, w_1190_, w_0896_);
xor (w_1905_, new_in1[1], new_in3[2]);
nand (w_1993_, w_0279_, w_1374_);
nand (w_1580_, w_1937_, w_1207_);
xor (w_1130_, new_in2[5], new_in4[1]);
or (w_0752_, w_2028_, w_1054_);
nand (w_0919_, w_0386_, w_1696_);
not (w_1228_, new_in10[3]);
nand (w_0960_, w_0947_, w_1460_);
nand (w_1235_, w_1713_, w_1096_);
nand (w_0554_, w_0691_, w_0584_);
nand (w_0792_, w_0527_, w_1826_);
xor (w_1683_, w_1381_, w_1995_);
nand (w_1908_, w_0348_, w_0764_);
nand (w_1829_, w_0863_, w_0886_);
and (w_0786_, w_1852_, w_1382_);
xor (w_1120_, w_1266_, w_2099_);
xor (w_0166_, new_in6[7], new_in3[2]);
xor (w_1046_, w_1931_, w_1904_);
nor (w_1114_, new_in10[2], new_in3[2]);
nand (w_1552_, w_1099_, w_0048_);
xor (w_0398_, w_1840_, w_0414_);
not (w_0352_, new_in9[3]);
nand (w_0164_, w_0726_, w_1051_);
nand (w_0869_, w_0200_, w_1535_);
xor (w_1540_, w_1930_, w_0571_);
and (w_1067_, new_in9[0], new_in1[0]);
and (w_1271_, w_1358_, w_1938_);
nand (w_1876_, w_1575_, w_0466_);
nand (w_1841_, w_0372_, w_1554_);
and (w_1837_, w_0225_, w_1298_);
nand (w_2036_, w_1545_, w_0338_);
xor (w_2032_, w_1411_, w_1463_);
xor (w_1501_, w_0636_, w_0387_);
nand (w_1887_, w_0018_, w_0345_);
nand (w_0709_, w_0485_, w_1501_);
nand (w_0521_, w_0596_, w_1247_);
nand (w_0971_, w_0035_, w_1762_);
or (w_0422_, w_0200_, w_0187_);
nand (w_0057_, w_0597_, w_0379_);
nand (w_0386_, new_in1[2], w_0333_);
nand (w_0615_, w_1708_, w_0191_);
nand (w_0604_, w_0168_, w_1592_);
nand (new_out3[1], w_1869_, w_0179_);
xor (w_0942_, w_0404_, w_2063_);
or (w_1996_, w_1860_, w_1935_);
nand (w_1674_, w_0605_, w_2030_);
nand (w_0406_, w_0168_, w_0898_);
nand (w_1549_, w_1707_, w_0420_);
and (w_0337_, new_in1[3], new_in3[1]);
xor (w_1083_, w_0381_, w_1627_);
and (w_1480_, w_0145_, w_2066_);
or (w_1278_, w_1243_, w_1510_);
nand (w_0305_, new_in1[1], new_in5[1]);
xor (w_1312_, w_0150_, w_1471_);
nand (w_1553_, w_1157_, w_1095_);
xor (w_0885_, new_in1[0], new_in3[3]);
nand (w_1871_, w_1708_, w_2035_);
xor (w_1342_, new_in5[7], new_in3[4]);
nand (w_1747_, w_0217_, w_0288_);
nand (w_2051_, w_1266_, w_2099_);
nand (w_2076_, w_0723_, w_1393_);
and (w_1599_, new_in11[0], new_in8[0]);
nand (w_0013_, w_1277_, w_0499_);
nor (w_1177_, new_in9[3], new_in1[0]);
and (w_0679_, new_in8[1], new_in9[4]);
and (w_0482_, w_1727_, w_1701_);
nand (w_1449_, w_0372_, w_0724_);
xor (w_0440_, w_0970_, w_0616_);
and (new_out1[2], w_0524_, w_0396_);
xor (w_0173_, w_2050_, new_in1[3]);
xor (w_1309_, new_in6[2], w_1165_);
xor (w_0583_, w_1198_, w_1512_);
xor (w_1191_, new_in2[6], new_in5[2]);
xor (w_2017_, new_in3[0], w_1001_);
xor (w_1736_, w_1112_, w_0330_);
nand (w_0182_, w_1860_, w_1935_);
xor (w_0140_, w_1706_, w_1743_);
nand (w_0012_, w_1734_, w_0988_);
xor (w_1660_, w_1228_, w_0062_);
and (w_1486_, w_0969_, w_1199_);
xor (w_1659_, w_0879_, w_1667_);
xor (w_0518_, w_0578_, w_0120_);
nand (w_0431_, w_1708_, w_0614_);
xor (w_1047_, new_in6[2], w_0745_);
xor (w_0707_, w_1716_, w_0946_);
nand (w_0131_, new_in8[3], w_1974_);
and (w_0263_, new_in10[0], new_in3[1]);
xor (w_0222_, w_0132_, w_1831_);
and (w_0239_, new_in10[1], new_in2[1]);
not (w_0580_, new_in2[0]);
xor (w_0365_, new_in4[3], new_in3[4]);
nand (w_0425_, w_0372_, w_0844_);
nand (w_1744_, w_0726_, w_1799_);
nand (w_2008_, w_0726_, w_0342_);
xor (w_1381_, new_in9[1], new_in1[1]);
and (w_1231_, w_0217_, w_1349_);
nand (w_0496_, w_1108_, w_0706_);
and (w_1375_, w_1527_, w_1409_);
xor (w_0710_, w_1259_, w_0622_);
xor (w_0540_, new_in9[1], new_in1[4]);
and (w_1204_, w_0052_, w_0994_);
xor (w_2053_, new_in6[1], w_1999_);
nand (w_0699_, w_0200_, w_1078_);
nand (w_0944_, w_0372_, w_1153_);
nand (w_0356_, w_0940_, w_1216_);
and (w_1431_, new_in10[1], new_in2[2]);
xor (w_1842_, new_in11[1], w_1511_);
nand (w_2000_, new_in3[0], w_2077_);
xor (w_1881_, w_2086_, w_0902_);
nand (w_0415_, w_0217_, w_0521_);
and (w_1020_, w_0721_, w_1376_);
nand (w_0106_, new_in6[3], w_0506_);
and (w_0943_, w_0217_, w_0564_);
and (new_out8[1], w_0922_, w_1906_);
xor (w_1057_, w_1848_, w_0542_);
nand (w_0084_, w_0200_, w_1229_);
xor (w_1936_, w_1767_, w_1342_);
xor (w_1978_, new_in6[8], new_in10[4]);
xor (w_1820_, w_0239_, w_0980_);
nand (w_1612_, w_1186_, w_1749_);
and (w_0082_, new_in9[1], new_in8[1]);
xor (w_0661_, new_in10[1], new_in7[1]);
and (new_out5[2], w_1367_, w_0504_);
or (w_1788_, w_1973_, w_0029_);
nand (w_0286_, new_in5[2], new_in2[3]);
or (w_0211_, new_in11[1], w_0100_);
nand (w_0019_, w_0058_, w_2049_);
xor (w_0074_, new_in5[1], new_in2[1]);
nand (w_0793_, w_0575_, w_2016_);
xor (w_0921_, w_0267_, w_0541_);
xor (w_0295_, w_1252_, new_in3[2]);
nand (w_1958_, new_in4[4], new_in10[4]);
xor (w_1586_, w_0876_, w_0076_);
nand (w_0015_, w_1354_, w_0884_);
xor (w_2090_, w_1350_, w_0568_);
nand (w_1386_, w_0578_, w_0120_);
nand (w_0989_, w_1699_, w_1640_);
xor (w_0750_, w_0360_, w_1637_);
xor (w_0808_, w_1879_, w_0737_);
and (w_1074_, w_0536_, w_1009_);
xor (w_1665_, w_1033_, w_1246_);
and (w_0314_, new_in6[1], new_in10[4]);
xor (w_0781_, new_in6[7], new_in2[2]);
xor (w_1831_, new_in11[1], new_in6[2]);
xor (w_1327_, w_0030_, w_0295_);
or (w_0027_, w_0200_, w_0203_);
xor (w_1827_, w_1061_, new_in5[4]);
nand (w_1303_, w_1796_, w_1094_);
nor (w_1108_, new_in6[1], new_in4[1]);
xor (w_2099_, new_in3[0], w_1129_);
or (w_1584_, w_0380_, w_1804_);
nand (w_0073_, w_1208_, w_0450_);
nand (w_1460_, w_1750_, w_0196_);
xor (w_0537_, w_0580_, w_0852_);
xor (w_0573_, w_1929_, w_0490_);
and (w_1214_, new_in6[2], new_in10[4]);
nand (w_1576_, w_0356_, w_1433_);
nand (w_0695_, w_1042_, new_in6[2]);
nand (w_1284_, w_1780_, w_1897_);
and (w_1060_, new_in4[0], w_0040_);
xor (w_1412_, w_1736_, w_0349_);
xor (w_0500_, w_1835_, w_1846_);
nor (w_0449_, w_0722_, w_1859_);
or (w_1893_, w_1833_, w_0668_);
nand (w_1112_, w_1519_, w_1351_);
xor (w_1879_, new_in6[1], new_in4[1]);
nand (w_0035_, w_0159_, w_1631_);
and (w_1149_, w_1784_, w_1497_);
nand (w_1757_, w_0200_, w_1829_);
xor (w_2063_, w_1946_, w_0730_);
nand (w_1170_, w_0586_, w_2003_);
nand (w_2029_, new_in6[1], new_in2[3]);
xor (w_0278_, w_1665_, w_0166_);
or (w_0618_, w_1375_, w_0139_);
xor (w_1755_, new_in9[2], new_in1[2]);
xor (w_1439_, w_0958_, w_0366_);
nand (w_0296_, w_1302_, w_1245_);
and (w_2085_, w_0983_, w_1492_);
xor (w_2089_, new_in4[5], w_0703_);
nand (w_0052_, new_in9[2], new_in1[5]);
nand (w_0857_, new_in1[0], w_1155_);
nand (w_0137_, w_0726_, w_0547_);
nand (w_0371_, w_0200_, w_0204_);
nor (w_1675_, new_in1[3], new_in9[6]);
xor (w_1885_, new_in1[1], new_in3[4]);
xor (w_1479_, w_0276_, w_2061_);
xor (w_1290_, new_in5[0], new_in2[4]);
or (w_1376_, w_1074_, w_0657_);
and (w_0741_, new_in5[1], new_in2[1]);
xor (w_0838_, new_in9[0], w_0312_);
xor (w_0283_, w_2097_, w_1455_);
xor (w_1706_, w_1003_, w_1430_);
or (w_1028_, w_0726_, w_2084_);
xor (w_0472_, new_in6[8], new_in3[3]);
nand (w_0213_, w_1427_, w_0719_);
xor (w_1818_, w_0487_, w_1255_);
nand (w_1692_, w_0716_, w_0791_);
nand (w_1437_, new_in8[3], new_in9[2]);
xor (w_1180_, new_in8[5], w_1377_);
or (w_1459_, w_1708_, w_2012_);
and (w_0442_, new_in3[0], new_in2[0]);
nand (w_1622_, w_0217_, w_1876_);
xor (w_2041_, w_0933_, w_1526_);
or (w_1068_, w_1913_, w_1110_);
nand (w_0115_, w_1841_, w_0577_);
nand (w_0998_, w_1593_, w_2059_);
xor (w_0797_, new_in6[5], new_in2[0]);
xor (w_0759_, new_in4[4], new_in1[2]);
xor (w_1811_, new_in10[2], w_1903_);
and (w_0349_, w_1942_, w_0437_);
nand (w_1094_, w_0984_, w_0689_);
and (w_1325_, new_in1[0], new_in8[5]);
and (w_1976_, new_in10[2], new_in4[2]);
xor (w_1615_, new_in10[0], new_in9[0]);
or (w_0149_, w_0954_, w_1855_);
nand (w_0293_, new_in2[2], new_in5[3]);
and (new_out7[3], w_0003_, w_1531_);
nand (w_0014_, w_1019_, w_1002_);
xor (w_1118_, w_1453_, w_1955_);
nand (w_1639_, w_2050_, new_in6[5]);
nand (w_0721_, w_1273_, w_1981_);
nand (w_0121_, new_in11[1], new_in7[1]);
and (w_1503_, new_in5[0], new_in2[0]);
xor (w_1955_, new_in6[2], new_in5[1]);
or (w_0575_, w_1879_, w_0006_);
not (w_1390_, w_0074_);
xor (w_1968_, w_0046_, w_0804_);
xor (w_0256_, w_1001_, w_1559_);
not (w_0336_, new_in5[8]);
xor (w_1276_, w_1254_, w_1405_);
and (w_1151_, w_1001_, w_1224_);
nand (w_0257_, w_0372_, w_1872_);
xor (w_1469_, new_in6[1], new_in2[5]);
and (w_0411_, w_1325_, w_0220_);
nand (w_0837_, w_0711_, w_1752_);
nand (w_0769_, w_2013_, w_0322_);
nand (w_0658_, w_0944_, w_0533_);
nand (w_0719_, w_1548_, w_0344_);
nand (w_0597_, w_0862_, w_2021_);
or (w_0530_, w_0726_, w_2090_);
and (w_2015_, w_0992_, w_1263_);
nand (w_0313_, w_1708_, w_0626_);
and (w_2028_, new_in5[2], new_in2[2]);
or (w_1772_, w_0726_, w_1026_);
xor (w_1321_, w_1253_, w_0601_);
xor (w_0641_, w_0967_, w_1515_);
xor (w_1542_, w_0123_, w_1577_);
nand (w_2075_, w_1708_, w_2074_);
xor (w_1126_, new_in2[5], new_in5[1]);
xor (w_1314_, w_0691_, w_0584_);
and (w_0277_, new_in10[0], w_0114_);
nand (w_1147_, new_in5[1], w_1560_);
nand (w_1556_, w_1056_, w_1352_);
nand (w_0056_, w_1505_, w_0553_);
xor (w_0049_, w_0599_, w_0620_);
xor (w_1132_, w_0357_, w_1027_);
nand (w_0549_, w_0200_, w_0704_);
or (w_1745_, w_0167_, w_0143_);
and (w_0951_, w_0954_, w_1441_);
nand (w_0455_, w_0252_, w_0518_);
not (w_1974_, new_in10[6]);
nand (w_0893_, new_in5[0], w_1928_);
nand (w_1059_, w_1595_, w_1929_);
nand (w_0531_, w_0717_, w_1150_);
nand (w_0515_, w_0200_, w_1359_);
and (w_0861_, new_in9[5], new_in8[0]);
xor (w_1730_, w_1887_, w_0473_);
nand (w_1316_, w_0092_, w_2045_);
nand (w_0591_, w_0678_, w_0710_);
nand (w_0810_, new_in2[5], new_in6[3]);
and (w_0433_, new_in3[3], new_in10[5]);
nand (w_1519_, new_in1[2], new_in3[2]);
xor (w_1502_, new_in3[3], w_2041_);
nand (w_0906_, new_in4[3], w_0258_);
nand (w_1257_, w_1211_, w_1132_);
xor (w_0973_, new_in8[2], new_in11[0]);
xor (w_0999_, new_in11[0], w_0701_);
and (w_1766_, w_0217_, w_0845_);
and (w_1550_, new_in8[3], new_in1[3]);
not (w_0513_, new_in2[5]);
nand (w_0147_, w_0200_, w_2015_);
nand (w_0266_, w_1665_, w_0166_);
nand (w_0065_, w_1878_, w_1102_);
or (w_1815_, w_1230_, w_0057_);
nand (w_1331_, w_1259_, w_0622_);
and (w_0471_, w_1379_, w_1657_);
not (w_1782_, new_in5[2]);
nand (w_0105_, w_1838_, w_0911_);
nand (w_0136_, new_in2[6], w_0932_);
nand (w_0933_, w_0497_, w_0229_);
xor (w_1505_, w_1833_, w_0668_);
nand (w_1878_, w_0726_, w_0816_);
nand (w_0638_, w_0726_, w_1394_);
xor (w_1626_, w_0976_, w_0608_);
and (w_1581_, new_in4[2], w_1165_);
and (w_1886_, w_0953_, w_1932_);
nand (w_1268_, w_1137_, w_1218_);
nand (w_0602_, w_1840_, w_0414_);
and (w_1203_, new_in10[4], new_in2[0]);
nor (w_2058_, w_2028_, w_1343_);
nand (w_1640_, w_1450_, w_0020_);
xor (w_0872_, new_in6[8], w_1960_);
nand (w_0694_, w_0372_, w_1057_);
xor (w_1154_, w_1296_, w_0359_);
nand (w_1942_, w_1929_, w_0490_);
nand (w_0434_, w_0168_, w_0465_);
nand (w_1701_, w_1832_, w_2056_);
nand (w_0637_, new_in10[1], new_in4[4]);
xor (w_1719_, w_0882_, w_1407_);
xor (w_1188_, w_0641_, w_1312_);
nand (w_0716_, w_1548_, w_0986_);
xor (w_0509_, w_0293_, w_1961_);
nand (w_1192_, new_in9[0], w_0312_);
and (w_1391_, w_1059_, w_0842_);
nand (w_0489_, new_in4[2], new_in3[3]);
or (w_1365_, w_1496_, w_1308_);
nand (w_0374_, w_0419_, w_1474_);
nand (w_2005_, w_2009_, w_1805_);
nand (w_0284_, w_0726_, w_0838_);
and (w_0090_, new_in8[0], w_0074_);
xor (w_0491_, w_0432_, w_1603_);
nand (w_0498_, w_0755_, new_in4[1]);
nand (w_1650_, new_in10[1], new_in3[4]);
xor (w_0894_, w_0846_, w_0058_);
or (w_1349_, w_0726_, w_0107_);
or (w_1596_, new_in4[3], w_0258_);
and (w_1765_, new_in10[3], new_in6[0]);
xor (w_0512_, new_in11[1], w_0080_);
nand (w_1251_, w_0200_, w_0786_);
xor (w_0830_, w_1983_, w_0685_);
xor (w_1894_, w_0925_, w_1408_);
xor (w_1027_, w_0058_, w_2049_);
nand (new_out6[0], w_0798_, w_0824_);
xor (w_1348_, new_in1[4], w_0629_);
xor (w_1498_, w_0800_, w_0424_);
nand (w_1176_, w_0821_, w_0346_);
and (w_0241_, w_1765_, w_1529_);
xor (w_0162_, w_0954_, w_1441_);
and (w_0550_, new_in8[4], new_in9[0]);
or (w_0022_, w_1513_, w_1953_);
xor (w_1293_, w_0951_, w_0500_);
xor (w_0187_, w_1894_, w_0945_);
nand (w_0232_, w_1708_, w_1475_);
nand (w_0897_, w_0735_, w_1340_);
nand (w_0647_, w_0200_, w_0854_);
nand (w_0497_, w_0367_, w_0891_);
nand (w_1854_, w_1480_, w_1726_);
xor (w_0478_, w_0775_, w_0242_);
nand (w_0678_, w_1723_, w_0709_);
xor (w_2055_, w_1557_, w_0797_);
nand (w_1593_, w_0726_, w_1116_);
or (w_0534_, w_1087_, w_1066_);
nand (w_0081_, w_1109_, w_0729_);
and (new_out5[1], w_0016_, w_1972_);
nand (w_0520_, w_1647_, w_0965_);
and (w_1105_, w_1645_, w_1284_);
and (w_0864_, new_in1[1], w_1598_);
and (w_1491_, w_0857_, w_1370_);
nand (w_1702_, w_1808_, w_2002_);
xor (w_0582_, w_0032_, w_0769_);
xor (w_1981_, w_1780_, w_1897_);
xor (w_0818_, w_1366_, w_1968_);
nand (w_0569_, w_1948_, w_0483_);
xor (w_2033_, w_0464_, w_0445_);
xor (w_0271_, new_in3[3], w_0795_);
xor (w_1789_, new_in10[4], w_1716_);
xor (w_0595_, new_in9[5], new_in8[5]);
and (w_1182_, w_1062_, w_0051_);
xor (w_2011_, new_in6[3], new_in4[3]);
not (w_0101_, w_0514_);
xor (w_0745_, w_1398_, w_0663_);
nor (w_1087_, w_1426_, w_1999_);
nand (w_1206_, w_0651_, w_1424_);
nand (w_1628_, w_0316_, w_0649_);
nand (w_1487_, w_0990_, w_0617_);
nand (w_0880_, new_in4[1], new_in5[5]);
and (w_0242_, w_1856_, w_0997_);
xor (w_1732_, w_1244_, w_0341_);
or (w_0186_, w_1509_, w_0593_);
and (w_0780_, w_1785_, w_0525_);
nand (w_1590_, w_0200_, w_1895_);
nand (w_0093_, w_0074_, w_1503_);
or (w_0778_, w_0123_, w_1073_);
xor (w_1055_, w_1647_, w_0965_);
nand (w_1926_, w_0623_, w_1616_);
xor (w_1474_, new_in1[1], new_in5[1]);
not (w_0030_, new_in10[5]);
nand (w_0048_, w_0726_, w_1710_);
nand (w_0174_, new_in1[2], new_in5[2]);
nand (w_1970_, w_0200_, w_2087_);
nand (w_0802_, new_in3[1], new_in2[1]);
nand (w_1152_, w_0503_, w_1303_);
nand (w_1752_, w_1883_, w_1686_);
nand (w_1708_, w_1965_, w_1774_);
nand (w_0731_, w_1797_, w_0548_);
nand (w_1261_, w_0201_, w_1329_);
xor (w_2038_, w_1212_, w_1055_);
nand (w_2056_, w_2039_, w_0894_);
xor (w_0917_, w_1406_, w_1730_);
xor (w_0867_, new_in3[3], w_1112_);
nand (w_1520_, w_2020_, w_0033_);
xor (w_0643_, w_0241_, w_0655_);
xor (w_0458_, w_0108_, w_0665_);
xor (w_1939_, w_1900_, w_1943_);
xor (w_1798_, w_0167_, w_0143_);
nand (new_out5[3], w_0422_, w_0549_);
xor (w_1259_, w_0326_, w_1423_);
xor (w_1687_, w_0566_, w_0949_);
xor (w_0982_, w_0040_, new_in5[4]);
xor (w_0223_, new_in2[3], new_in7[0]);
nand (w_0974_, w_0315_, w_0887_);
or (w_1852_, w_1708_, w_0475_);
nand (w_0791_, w_0726_, w_1901_);
xor (w_0588_, w_0189_, w_1842_);
nand (w_0722_, w_2036_, w_0476_);
xor (w_0462_, w_1926_, w_0645_);
and (w_1007_, w_1835_, w_1846_);
xor (w_1029_, w_0063_, w_0472_);
not (w_1273_, w_1929_);
nand (w_1270_, w_0186_, w_1672_);
xor (w_0936_, w_2027_, w_1633_);
xor (w_1004_, w_1163_, w_0393_);
nand (w_1127_, w_1548_, w_1014_);
xor (w_0825_, w_0040_, new_in5[3]);
xor (w_0420_, w_0741_, w_1373_);
or (w_1208_, w_0217_, w_1439_);
nand (w_0798_, w_0200_, w_0733_);
and (w_2062_, w_1459_, w_0206_);
nand (w_0129_, w_1362_, w_1436_);
nand (new_out10[1], w_1494_, w_0176_);
nand (w_0053_, w_1857_, w_0224_);
xor (w_1716_, new_in8[1], new_in3[1]);
and (w_0868_, w_1525_, w_1611_);
and (w_0795_, new_in4[7], new_in10[4]);
xor (w_0123_, new_in2[6], new_in5[7]);
and (w_1602_, w_0217_, w_0409_);
xor (w_1691_, w_0388_, w_0184_);
xor (w_1690_, new_in6[4], w_0106_);
or (w_1685_, new_in1[1], new_in9[4]);
or (w_1699_, w_0217_, w_1065_);
xor (w_1751_, w_1719_, w_0274_);
nand (w_0170_, w_0726_, w_0606_);
nand (w_1769_, new_in11[1], w_0080_);
and (w_1997_, new_in4[5], new_in10[2]);
and (w_1558_, w_1235_, w_0779_);
nand (w_0966_, w_0241_, w_0655_);
xor (w_0237_, w_1232_, w_0867_);
nand (w_1402_, w_0168_, w_0156_);
and (w_0054_, new_in5[0], w_1885_);
xor (w_0417_, w_1939_, w_0750_);
nand (w_0623_, w_0920_, w_1798_);
nand (w_0723_, w_0768_, w_0924_);
nand (w_1239_, w_0442_, w_0562_);
xor (w_0490_, w_0023_, w_1250_);
and (w_0168_, w_1123_, w_1270_);
xor (w_1077_, w_1539_, w_1811_);
nand (w_0782_, w_1288_, w_0895_);
nand (w_1364_, new_in4[3], new_in1[1]);
xor (w_0366_, w_1324_, w_0753_);
nand (w_0610_, w_0217_, w_1989_);
xor (w_0461_, w_2042_, w_1015_);
nand (w_1525_, w_1815_, w_1486_);
and (w_1410_, w_1256_, w_0615_);
and (w_0511_, new_in3[0], new_in2[1]);
or (w_1340_, new_in2[5], new_in6[3]);
nand (w_0711_, new_in9[3], new_in1[2]);
xor (w_0611_, w_0446_, w_0968_);
and (w_0446_, w_1437_, w_1152_);
and (w_1243_, w_0136_, w_0742_);
xor (w_1792_, new_in4[0], w_0783_);
xor (w_0608_, new_in9[3], w_1293_);
xor (w_0058_, new_in5[1], new_in2[2]);
xor (w_0438_, new_in11[0], new_in8[0]);
nand (w_1808_, w_1022_, w_1912_);
xor (w_0224_, new_in7[0], w_1881_);
not (w_1630_, new_in10[2]);
nand (w_0350_, new_in6[1], new_in4[1]);
nand (w_0159_, w_0706_, w_0134_);
nor (w_1049_, w_0888_, w_1332_);
xor (w_1582_, new_in1[3], new_in3[3]);
nand (w_1680_, w_0217_, w_1993_);
or (w_0969_, w_0935_, w_1721_);
nand (w_1428_, w_0372_, w_1676_);
xor (w_1929_, w_0149_, w_2081_);
and (w_0155_, new_in6[0], new_in10[6]);
or (w_1880_, w_0613_, w_0833_);
xor (w_0362_, w_1561_, w_1315_);
xor (w_1397_, w_1877_, w_0528_);
not (w_1693_, new_in4[7]);
or (w_1836_, w_0726_, w_2007_);
xor (w_1467_, new_in4[0], new_in5[4]);
nand (w_0803_, w_1925_, new_in1[1]);
or (w_0018_, w_0046_, w_0804_);
and (w_1767_, new_in3[3], new_in5[6]);
xor (w_0762_, new_in9[2], new_in1[0]);
nand (w_0046_, w_0538_, w_0255_);
xor (w_0548_, w_0492_, w_1222_);
nand (w_0190_, w_0403_, w_0682_);
xor (w_0165_, new_in5[1], new_in6[5]);
nand (w_1698_, w_1472_, w_2019_);
nand (w_0436_, w_1857_, w_0916_);
nand (w_1507_, w_0598_, w_0028_);
xor (w_1695_, w_1828_, w_2077_);
not (w_0430_, w_0531_);
and (w_1110_, w_0205_, w_0720_);
xor (w_0370_, w_1862_, w_0866_);
xor (w_0113_, w_0827_, w_1417_);
and (w_0195_, w_0077_, w_1420_);
nand (w_0483_, w_0217_, w_1770_);
xor (w_1888_, new_in8[4], w_0480_);
or (w_0585_, w_0862_, w_1923_);
and (w_0357_, w_0393_, w_1045_);
xor (w_0388_, w_1052_, w_0058_);
nand (w_1450_, w_1548_, w_1134_);
nand (w_1353_, new_in11[1], new_in6[2]);
nand (w_0673_, w_0168_, w_1258_);
or (w_0145_, new_in9[0], new_in8[0]);
nand (w_1462_, new_in2[6], new_in5[7]);
and (w_1117_, new_in6[2], w_1165_);
nand (w_0599_, w_1008_, w_1617_);
nand (w_0310_, w_1681_, w_0624_);
nand (w_0596_, w_1548_, w_0659_);
and (w_1839_, new_in3[1], w_1997_);
xor (w_0243_, w_1685_, w_1490_);
xor (w_0407_, new_in3[2], w_0788_);
nand (w_2079_, w_1708_, w_2070_);
xor (w_1339_, w_0676_, w_1048_);
xor (w_1070_, w_0789_, w_0207_);
nand (w_1534_, w_2096_, w_0808_);
nand (w_0033_, w_1548_, w_0194_);
xor (w_1495_, w_0613_, w_0833_);
xor (w_1509_, w_2085_, w_1555_);
and (w_1000_, new_in8[4], new_in9[1]);
xor (w_1254_, w_0771_, w_0429_);
xor (w_0544_, w_0467_, w_1435_);
xor (w_0923_, w_0068_, w_0523_);
nand (w_1351_, w_0149_, w_2081_);
nand (w_0346_, w_0056_, w_0081_);
xor (w_0460_, new_in3[4], w_0478_);
xor (w_0156_, w_0678_, w_0710_);
xor (w_1202_, w_0507_, w_1783_);
nand (w_1341_, w_1708_, w_1395_);
xor (w_0965_, w_1913_, w_1689_);
xor (w_0292_, w_0706_, w_0134_);
xor (w_1892_, w_0090_, w_2037_);
or (w_0832_, w_0447_, w_1986_);
nand (w_1579_, w_1857_, w_0171_);
nand (w_1954_, w_0200_, w_1724_);
not (w_2050_, new_in4[5]);
nand (w_1414_, w_1698_, w_0278_);
nand (w_0358_, w_0372_, w_1664_);
nand (w_1648_, w_0880_, w_2094_);
nand (w_0282_, w_0726_, w_1963_);
nand (w_0212_, w_2005_, w_0009_);
nand (w_1267_, w_1716_, w_0946_);
nand (w_0070_, new_in2[4], new_in5[2]);
nand (w_1623_, new_in3[1], w_1148_);
and (w_0096_, new_in9[4], new_in8[0]);
xor (w_0157_, w_1432_, w_0043_);
xor (w_0785_, w_0993_, w_2068_);
nand (w_0994_, w_0531_, w_1758_);
xor (w_0249_, w_1469_, w_1615_);
xor (w_1383_, w_2067_, w_0981_);
xor (w_1889_, new_in10[1], new_in3[4]);
and (w_1289_, new_in8[4], new_in1[0]);
and (w_0836_, new_in5[0], new_in5[1]);
nand (w_0427_, w_1422_, w_1024_);
or (w_0903_, w_1545_, w_0010_);
and (w_0811_, w_0495_, w_0153_);
xor (w_0654_, w_0503_, w_1303_);
and (w_0625_, w_2052_, w_0309_);
and (w_1689_, new_in5[1], new_in2[2]);
xor (w_0851_, w_1452_, w_1111_);
or (w_0177_, w_0046_, w_0244_);
xor (w_0995_, new_in5[1], new_in5[2]);
nand (w_0148_, w_0827_, new_in9[2]);
xor (w_1357_, w_0560_, w_0169_);
or (w_1657_, w_1013_, w_1092_);
and (w_0840_, w_0199_, w_1547_);
xor (w_1758_, new_in9[2], new_in1[5]);
or (w_0039_, w_1345_, w_0900_);
nand (w_0747_, w_1857_, w_0936_);
xor (w_0688_, new_in6[4], new_in4[8]);
nand (w_1446_, w_1778_, w_0930_);
nand (w_1297_, new_in6[6], new_in7[1]);
or (w_0051_, w_1034_, w_0805_);
not (w_0368_, w_1300_);
xor (w_0028_, w_1000_, w_0928_);
xor (w_2086_, new_in3[0], new_in2[0]);
nand (w_1477_, w_1361_, w_1363_);
nand (w_1807_, w_0200_, w_1039_);
nand (w_1358_, w_1431_, w_1160_);
xor (w_2066_, new_in5[0], new_in2[0]);
xor (w_1456_, w_0920_, w_1798_);
nand (w_0896_, w_1708_, w_1908_);
and (w_0384_, new_in6[1], w_0513_);
and (w_1345_, w_0070_, w_1347_);
xor (w_1423_, w_0129_, w_1191_);
xor (w_0193_, new_in4[1], new_in5[5]);
not (w_1921_, new_in6[1]);
xor (w_1144_, w_2039_, w_0894_);
nor (w_1714_, w_0185_, w_0511_);
nand (w_0328_, w_1084_, w_0170_);
and (w_1107_, new_in10[2], new_in2[2]);
xor (w_1949_, new_in8[1], w_0435_);
and (w_2059_, w_0217_, w_1532_);
and (w_0238_, new_in5[1], new_in2[3]);
xor (w_0456_, new_in11[1], w_1498_);
nand (new_out10[2], w_1759_, w_1402_);
and (w_0325_, new_in1[1], new_in3[2]);
xor (w_0260_, w_0046_, w_0707_);
xor (w_0834_, new_in9[3], new_in1[3]);
nand (w_1076_, w_0901_, w_1333_);
nand (w_1041_, w_0739_, w_1240_);
nand (w_1786_, w_0217_, w_1299_);
nand (w_1663_, w_0007_, w_0754_);
xor (w_0272_, w_1600_, w_0353_);
xor (w_0657_, w_1929_, w_1981_);
and (w_1301_, w_0552_, w_1488_);
xor (w_0634_, new_in10[1], new_in6[5]);
and (w_1875_, w_1158_, w_0148_);
or (w_1002_, w_0901_, w_1333_);
and (w_1577_, w_0484_, w_0585_);
xor (w_1966_, w_0827_, w_0079_);
and (w_0285_, w_1596_, w_2073_);
xor (w_0475_, w_0075_, w_1215_);
nand (w_2078_, w_0741_, w_1113_);
xor (w_1095_, new_in6[2], w_1337_);
xor (w_0333_, w_1087_, w_1066_);
nand (w_0441_, w_0168_, w_0914_);
or (w_0516_, w_1060_, w_1130_);
xor (w_1735_, w_1345_, w_0900_);
xor (w_1511_, w_0644_, w_1683_);
nor (w_0185_, new_in3[0], new_in2[1]);
or (w_1717_, w_1649_, w_1602_);
and (w_1835_, new_in1[0], new_in3[3]);
xor (w_1741_, w_1056_, w_1352_);
nand (w_0651_, w_0217_, w_0687_);
xor (w_1709_, w_1397_, w_1182_);
xor (w_0701_, w_1503_, w_0634_);
nand (w_0819_, w_0372_, w_1691_);
xor (w_1017_, new_in2[1], w_0410_);
nand (w_1445_, w_0357_, w_1027_);
xor (w_1442_, w_1108_, w_0706_);
nand (w_0627_, w_0142_, w_1399_);
xor (w_0245_, w_0347_, w_0573_);
and (w_1064_, new_in6[0], new_in10[4]);
nand (w_0718_, w_1708_, w_1565_);
nand (w_1295_, w_1306_, w_0329_);
and (w_0220_, new_in8[4], new_in1[1]);
nand (w_0705_, new_in4[0], new_in1[2]);
xor (w_1136_, new_in6[7], new_in5[3]);
xor (w_1443_, new_in10[0], w_2053_);
nand (w_0815_, w_1297_, w_1663_);
nand (w_0809_, w_0832_, w_1748_);
and (w_0656_, w_1174_, w_0314_);
nand (w_0299_, w_0302_, w_0428_);
xor (w_0831_, w_1833_, w_0433_);
not (w_0488_, new_in4[6]);
xor (w_0207_, new_in4[4], new_in10[4]);
and (w_0311_, w_0662_, w_0294_);
xor (w_0203_, w_1765_, w_1529_);
nor (w_1260_, w_0205_, w_0720_);
nand (w_0178_, w_1212_, w_1055_);
and (w_1613_, new_in4[0], new_in8[0]);
nand (w_0279_, w_0726_, w_0766_);
xor (w_0029_, new_in10[2], new_in9[4]);
xor (w_1633_, new_in10[0], new_in4[0]);
xor (w_0579_, new_in9[4], new_in1[3]);
nand (w_0779_, w_1725_, w_1891_);
nand (w_0341_, w_0539_, w_1612_);
xor (w_0042_, new_in3[2], new_in2[3]);
xor (w_2084_, w_1977_, w_1874_);
xor (w_1346_, new_in1[2], w_0333_);
nor (w_1315_, w_1976_, w_0031_);
nand (w_0768_, w_1936_, w_1820_);
and (w_0276_, w_0958_, w_1244_);
nand (w_0653_, w_0168_, w_1746_);
nand (new_out3[2], w_1106_, w_0660_);
nand (w_0905_, w_0310_, w_1193_);
xor (w_0382_, new_in3[3], new_in5[6]);
xor (w_1661_, w_0723_, w_1393_);
nor (w_1931_, w_0987_, w_1810_);
nand (w_1863_, w_1969_, w_0451_);
or (w_1044_, w_1572_, w_1625_);
or (w_1715_, w_0217_, w_0185_);
and (w_0551_, w_1462_, w_0501_);
xor (w_1986_, w_1137_, w_1221_);
nand (w_1361_, new_in11[1], w_1498_);
nand (w_1185_, w_1295_, w_1248_);
and (w_0823_, w_2086_, w_0902_);
and (w_1359_, w_1914_, w_0927_);
nand (w_1694_, w_1708_, w_1365_);
nand (w_1418_, w_0823_, w_1118_);
xor (w_1605_, w_1684_, w_0452_);
nand (w_0198_, w_1708_, w_1388_);
xor (w_1368_, w_0270_, w_1017_);
nand (w_2093_, w_1213_, w_1788_);
and (w_0945_, w_1551_, w_1281_);
xor (w_0034_, w_2001_, w_1456_);
nand (w_0180_, new_in6[3], w_0862_);
and (w_0835_, w_0217_, w_1564_);
xor (w_0494_, new_in10[4], new_in7[1]);
xor (w_1515_, new_in6[4], new_in2[8]);
nand (w_1538_, w_0251_, w_0796_);
xor (w_0235_, new_in6[2], new_in2[4]);
xor (w_1167_, new_in10[1], new_in9[1]);
and (w_1629_, new_in8[3], new_in1[1]);
and (w_0404_, w_1170_, w_1482_);
and (w_0354_, new_in5[0], new_in2[4]);
xor (w_1991_, w_0522_, w_1421_);
nand (w_0229_, w_1225_, w_1793_);
nand (w_1979_, new_in9[4], new_in1[3]);
xor (w_0631_, new_in9[6], new_in8[6]);
and (w_1217_, new_in11[0], w_0352_);
and (w_1928_, new_in5[1], w_1782_);
xor (w_0866_, w_0586_, w_2003_);
and (w_1052_, new_in5[0], new_in2[1]);
xor (w_0273_, w_1646_, w_1761_);
nand (w_0739_, new_in2[6], new_in5[2]);
nand (w_0635_, w_1548_, w_1083_);
xor (w_0663_, new_in10[1], w_1542_);
nand (w_1135_, w_0200_, w_0658_);
xor (w_1667_, new_in2[6], new_in4[2]);
xor (w_0881_, new_in9[5], new_in1[2]);
nand (w_0970_, w_1802_, w_0777_);
nand (w_0794_, w_0299_, w_1136_);
and (w_1523_, w_0702_, w_0382_);
and (w_1216_, new_in5[8], w_1069_);
nand (w_0744_, w_0728_, w_2043_);
not (w_1925_, new_in9[1]);
or (w_1248_, w_1306_, w_0329_);
nand (w_1237_, w_1857_, w_2082_);
xor (w_0381_, new_in9[0], new_in8[1]);
or (w_0439_, new_in11[1], w_0010_);
and (w_0167_, new_in10[0], w_0529_);
and (w_0784_, new_in8[2], new_in9[2]);
xor (w_0002_, w_0715_, w_1334_);
and (w_0713_, new_in10[0], new_in3[3]);
nand (w_0418_, w_1693_, new_in6[3]);
nand (w_1864_, w_0376_, w_1144_);
nand (w_0626_, w_1058_, w_1316_);
xor (w_2068_, new_in8[0], new_in7[0]);
xor (w_1011_, w_0026_, w_0122_);
xor (w_1826_, new_in4[0], w_1326_);
or (w_1567_, w_1435_, w_1114_);
xor (w_1153_, w_1249_, w_0666_);
xor (w_0355_, w_0813_, w_0680_);
and (w_1209_, w_1913_, w_1689_);
nand (w_1198_, w_1257_, w_0296_);
or (w_1932_, w_0026_, w_0122_);
nand (w_1146_, new_in8[3], new_in9[3]);
xor (w_0527_, w_0430_, w_1758_);
and (w_0796_, w_0217_, w_0282_);
or (w_1264_, w_1689_, w_0078_);
xor (w_0895_, w_0861_, w_0679_);
xor (w_0104_, w_1910_, w_1030_);
or (w_0742_, w_0384_, w_0304_);
xor (w_1592_, w_0237_, w_1391_);
and (w_0743_, w_1028_, w_0736_);
xor (w_1448_, new_in8[6], w_1305_);
or (w_0390_, w_0689_, w_1917_);
nand (w_1722_, w_1068_, w_0226_);
xor (w_1506_, w_1480_, w_1726_);
nand (w_1773_, w_1280_, w_1413_);
and (w_0059_, new_in1[0], new_in3[4]);
xor (w_0320_, new_in3[4], new_in1[4]);
xor (w_0143_, new_in10[1], new_in9[3]);
nand (w_0303_, w_0217_, w_1543_);
xor (w_1134_, w_1729_, w_0772_);
xor (w_1245_, w_1211_, w_1132_);
or (w_0448_, w_1797_, w_0548_);
nand (w_1585_, new_in6[7], new_in5[3]);
nand (w_1461_, w_1401_, w_0526_);
xor (w_1258_, new_in10[2], new_in4[1]);
xor (w_1676_, w_0438_, w_0165_);
xor (w_1655_, w_0527_, w_1826_);
nand (w_0983_, w_1693_, new_in6[7]);
xor (w_0004_, new_in2[6], new_in6[4]);
or (w_0961_, w_1337_, w_0408_);
nand (w_1106_, w_0200_, w_0197_);
nand (w_1642_, w_0372_, w_1763_);
nand (w_0088_, new_in8[1], new_in11[1]);
nand (w_1677_, new_in9[5], w_0878_);
or (w_0841_, w_1546_, w_0909_);
nand (w_1614_, w_0054_, w_0124_);
xor (w_1215_, new_in4[0], new_in3[1]);
and (w_0928_, new_in9[0], new_in8[5]);
or (w_0758_, w_0726_, w_1412_);
xor (w_1935_, w_1863_, w_1518_);
xor (w_1012_, w_1166_, w_1756_);
not (w_1161_, new_in10[1]);
xor (w_1091_, w_0973_, w_0762_);
nand (w_1819_, w_1483_, w_1169_);
not (w_1545_, new_in11[1]);
xor (w_1524_, w_1074_, w_0657_);
nand (w_1578_, w_1449_, w_0592_);
xor (w_0848_, w_0263_, w_1884_);
xor (w_2046_, w_0046_, w_1588_);
nand (w_0339_, w_0168_, w_1951_);
nand (w_0024_, w_1708_, w_0667_);
nand (w_0930_, w_1419_, w_1843_);
nand (w_0506_, w_1353_, w_0570_);
and (w_1219_, w_1386_, w_0455_);
nand (w_0045_, w_1127_, w_0943_);
or (w_0729_, w_1505_, w_0553_);
nand (w_2087_, w_0890_, w_1090_);
nand (w_0288_, w_0373_, w_1400_);
nand (w_0570_, w_0132_, w_1831_);
nand (w_2088_, new_in8[1], w_0706_);
nand (w_1933_, w_1545_, w_1511_);
nand (w_1738_, w_1896_, w_0807_);
and (w_1229_, w_1624_, w_0313_);
nand (w_0302_, new_in6[6], new_in5[2]);
nand (w_0291_, w_1089_, w_1918_);
nand (w_0199_, w_0827_, new_in10[6]);
xor (w_0632_, new_in8[3], w_2017_);
xor (w_1961_, w_0286_, w_0767_);
and (w_2042_, w_0951_, w_0500_);
nand (w_1631_, w_1283_, w_0292_);
nand (w_1938_, w_1195_, w_0038_);
nand (w_1869_, w_0200_, w_0280_);
xor (w_0909_, new_in4[5], new_in6[5]);
xor (w_1746_, w_0443_, w_1470_);
xor (w_0562_, new_in3[1], new_in2[1]);
or (w_1162_, w_0217_, w_0130_);
and (w_2045_, w_0217_, w_0137_);
xor (w_0666_, w_0243_, w_0046_);
xor (w_0219_, w_0609_, w_0111_);
xor (w_0828_, w_1875_, w_1845_);
and (w_1883_, new_in9[2], new_in1[1]);
xor (w_0968_, w_0013_, w_0683_);
nand (w_1432_, w_1643_, w_0684_);
nand (w_0423_, w_0200_, w_1410_);
xor (w_0720_, new_in5[2], new_in2[1]);
not (w_0372_, w_1708_);
nand (w_0196_, w_1608_, w_1467_);
xor (w_0269_, w_0594_, w_1544_);
nand (w_2073_, new_in6[3], w_0906_);
and (w_1743_, w_0671_, w_2076_);
nand (w_0664_, w_1115_, w_0748_);
nand (w_0536_, w_1287_, w_2038_);
nand (w_1748_, w_0731_, w_0363_);
nand (w_1725_, w_0908_, w_1418_);
xor (w_1891_, w_1713_, w_1096_);
nand (w_1433_, w_1076_, w_0014_);
and (w_0132_, new_in6[1], new_in11[0]);
and (w_0737_, new_in10[4], new_in3[2]);
nand (w_1959_, w_0726_, w_0561_);
xor (w_1015_, w_1007_, w_0746_);
and (w_1003_, w_0873_, w_1702_);
nand (w_0450_, w_0217_, w_1520_);
nand (w_1016_, w_1958_, w_0849_);
or (w_1742_, w_1679_, w_0937_);
xor (w_1601_, w_0650_, w_1732_);
or (w_0975_, w_0217_, w_0557_);
nand (w_0044_, w_0467_, w_1435_);
xor (w_0568_, new_in5[0], new_in1[0]);
and (w_1140_, w_0217_, w_0874_);
nor (w_1784_, w_0595_, w_0633_);
xor (w_0732_, w_0556_, w_0444_);
nand (w_0221_, w_2094_, w_1043_);
xor (w_0234_, new_in8[5], w_0405_);
nand (w_0373_, w_1548_, w_0083_);
nand (w_1724_, w_0672_, w_1844_);
xor (w_0929_, w_1384_, w_1203_);
nand (w_1822_, w_0005_, w_0236_);
nand (w_1707_, new_in8[4], new_in4[6]);
xor (w_1999_, new_in2[3], new_in5[4]);
and (w_1225_, w_1469_, w_1615_);
nand (w_0077_, w_0827_, w_0459_);
xor (w_0727_, new_in6[8], new_in5[4]);
nand (w_1800_, new_in11[1], w_0100_);
nand (new_out3[0], w_1175_, w_0339_);
nand (w_1197_, w_1857_, w_0460_);
nand (w_0385_, new_in8[1], w_1373_);
not (w_0075_, new_in8[0]);
xor (w_0561_, w_1067_, w_1975_);
and (w_1828_, new_in10[2], new_in4[1]);
nand (w_1564_, w_0102_, w_2008_);
xor (w_1111_, w_1220_, w_1589_);
xor (w_1466_, w_1325_, w_0220_);
xor (w_0555_, w_0411_, w_1276_);
nand (w_1522_, w_1857_, w_0064_);
nand (w_1809_, w_0168_, w_1188_);
xor (w_0644_, w_0463_, w_1635_);
and (w_0078_, w_1052_, w_0058_);
and (w_0258_, w_0695_, w_1893_);
nand (w_1150_, w_0751_, w_0540_);
xor (w_0993_, w_0114_, new_in1[0]);
nand (w_1299_, w_0758_, w_0532_);
nand (w_1597_, new_in10[1], new_in7[1]);
xor (w_0445_, w_1974_, w_2044_);
xor (w_0914_, w_1098_, w_1660_);
xor (w_0681_, new_in10[2], new_in9[2]);
or (w_2083_, w_1708_, w_0926_);
nand (w_1956_, w_1440_, w_0530_);
xor (w_1010_, w_1177_, w_2023_);
xor (w_1500_, w_0529_, w_0273_);
xor (w_0714_, w_0075_, new_in3[0]);
xor (w_0240_, w_1138_, w_0509_);
xor (w_1096_, new_in6[3], new_in5[2]);
xor (w_1666_, new_in9[4], w_0461_);
nand (w_1210_, new_in4[2], new_in5[6]);
xor (w_0941_, new_in5[0], w_1885_);
xor (w_1403_, w_1973_, w_0029_);
or (w_1624_, w_1708_, w_0588_);
xor (w_0612_, w_0755_, new_in5[3]);
and (w_1669_, new_in10[3], new_in6[1]);
xor (w_1453_, w_0442_, w_0562_);
nand (w_1422_, w_0372_, w_0581_);
nand (new_out7[2], w_0371_, w_1223_);
nor (w_2034_, new_in8[3], new_in9[3]);
nand (w_0248_, w_0381_, w_1627_);
nand (w_0287_, new_in10[1], new_in3[2]);
nand (w_0687_, w_1200_, w_0098_);
xor (w_0628_, w_1186_, w_1749_);
xor (w_0991_, w_1678_, w_1754_);
xor (w_1705_, w_0545_, w_0285_);
nand (w_0662_, new_in2[5], new_in5[6]);
nand (w_1452_, w_0468_, w_1940_);
or (w_0160_, w_0217_, w_1476_);
xor (w_0447_, w_0735_, w_0642_);
xor (w_0986_, w_1795_, w_0512_);
and (w_1272_, w_1567_, w_1571_);
and (w_0962_, w_1644_, w_0830_);
nand (w_1565_, w_0648_, w_0619_);
nand (w_0574_, w_1708_, w_0474_);
nand (w_0389_, w_1143_, w_0135_);
xor (w_1504_, w_1673_, w_1404_);
xor (w_1336_, new_in10[3], new_in4[3]);
or (w_0412_, w_0726_, w_0066_);
nand (w_0875_, w_1548_, w_0603_);
xor (w_1006_, new_in8[3], new_in11[1]);
xor (w_1404_, w_0082_, w_0355_);
nand (w_0814_, w_1708_, w_0989_);
xor (w_1951_, w_0958_, w_1244_);
nand (w_2009_, w_1719_, w_0274_);
nand (w_0468_, w_1310_, w_1403_);
and (w_1734_, new_in4[0], new_in3[1]);
and (w_1398_, new_in10[0], w_1447_);
xor (w_0542_, w_0827_, w_1740_);
nand (w_0860_, w_0200_, w_1578_);
and (w_1913_, new_in5[2], new_in2[1]);
nand (w_0749_, w_0036_, w_1641_);
nand (w_1753_, new_in4[4], new_in1[2]);
nand (w_1604_, w_1688_, w_0910_);
xor (w_0636_, w_1050_, w_0172_);
nand (w_1616_, w_2001_, w_1456_);
and (w_1644_, w_1669_, w_1064_);
and (w_1806_, w_1331_, w_0591_);
and (w_0948_, w_1812_, w_0820_);
or (w_1420_, w_1651_, w_1415_);
xor (w_1171_, w_1674_, w_0544_);
nand (w_0069_, w_0182_, w_0868_);
or (w_0790_, w_1708_, w_1605_);
xor (w_0902_, new_in5[0], new_in6[1]);
xor (w_0775_, w_0641_, w_0049_);
nand (w_0947_, w_0301_, w_0221_);
nand (w_1847_, w_0418_, w_0618_);
nand (w_1131_, new_in10[2], new_in3[5]);
and (new_out11[3], w_0200_, w_0015_);
nand (w_1380_, w_1857_, w_0942_);
nand (w_1274_, w_0200_, w_1294_);
nand (w_0154_, w_1909_, w_1944_);
nand (w_1371_, w_0343_, w_2025_);
nand (w_1137_, w_1210_, w_0996_);
nand (w_0884_, w_1708_, w_1371_);
nand (w_1830_, w_0976_, w_0608_);
and (w_1791_, w_1131_, w_1196_);
nand (w_1298_, w_0372_, w_1670_);
nand (w_1175_, w_0200_, w_1919_);
xor (w_0502_, w_0138_, w_1282_);
or (w_0912_, w_0621_, w_1500_);
nand (w_1249_, w_1010_, w_1001_);
nand (w_0201_, new_in8[2], new_in4[2]);
and (w_1740_, new_in8[2], w_1227_);
xor (w_1526_, w_0395_, w_0477_);
xor (w_2002_, new_in5[8], new_in3[5]);
xor (w_0547_, w_0109_, w_1751_);
xor (w_0443_, w_0326_, w_1368_);
xor (w_0546_, new_in7[1], w_0799_);
or (w_0476_, w_1217_, w_0188_);
nand (w_1277_, new_in4[3], new_in10[4]);
xor (w_1678_, w_0036_, w_1978_);
xor (w_0624_, new_in1[2], new_in3[3]);
nand (w_1189_, w_0904_, w_0793_);
and (w_0094_, w_0489_, w_0664_);
nand (w_2071_, w_0372_, w_0458_);
nand (w_0767_, new_in2[4], new_in5[1]);
xor (w_1529_, w_1001_, w_0393_);
nand (w_0192_, w_0670_, w_1766_);
nand (w_0859_, w_0168_, w_1320_);
nand (w_1213_, w_1630_, new_in9[4]);
nand (w_1201_, new_in4[1], new_in3[2]);
or (w_0504_, w_0200_, w_1731_);
and (w_1952_, w_1983_, w_0685_);
xor (w_0080_, w_1651_, w_1415_);
nand (w_0011_, w_0713_, w_1889_);
xor (w_1635_, new_in8[1], new_in7[1]);
nand (w_0646_, w_0800_, w_0424_);
nand (w_1851_, w_0639_, w_0635_);
not (w_1061_, new_in2[3]);
and (w_0426_, w_2069_, w_1994_);
and (w_1774_, w_0216_, w_0840_);
nand (w_0953_, w_1434_, w_0219_);
xor (w_0958_, new_in1[0], new_in3[0]);
xor (w_1963_, w_1117_, w_0140_);
nand (w_0003_, w_0200_, w_1837_);
xor (w_0009_, w_0843_, w_0261_);
and (w_0858_, new_in9[0], new_in8[6]);
nand (w_0008_, w_1900_, w_1943_);
nand (w_0849_, w_0789_, w_0207_);
and (w_1103_, new_in4[0], new_in5[4]);
xor (w_0095_, w_0598_, w_0028_);
nand (w_0421_, new_in8[2], new_in3[2]);
and (w_1917_, w_0114_, new_in8[1]);
nand (w_2020_, w_0726_, w_0001_);
nand (w_2021_, w_0514_, w_0025_);
xor (w_1490_, w_0713_, w_1889_);
nand (w_0855_, w_0360_, w_1637_);
xor (w_1861_, w_1755_, w_1082_);
or (w_0060_, w_1925_, w_0260_);
nand (w_1912_, w_1767_, w_1342_);
nand (w_0191_, w_0394_, w_1292_);
nand (w_2069_, new_in3[2], w_0788_);
nand (w_1081_, w_1337_, w_0408_);
xor (w_1093_, w_1225_, w_1793_);
xor (w_0799_, w_0823_, w_1118_);
xor (w_0454_, w_0956_, w_0761_);
xor (w_1603_, new_in1[3], w_0972_);
xor (w_1760_, w_1159_, w_1813_);
xor (w_1943_, new_in8[1], w_0706_);
xor (w_1378_, w_0929_, w_1271_);
or (w_1834_, w_1280_, w_1413_);
xor (w_1045_, new_in6[1], new_in4[5]);
xor (w_0103_, w_1013_, w_1092_);
xor (w_1030_, w_0555_, w_1550_);
nand (w_1899_, w_1879_, w_1810_);
and (w_0801_, new_in2[1], new_in5[4]);
xor (w_0692_, w_1473_, w_1654_);
nand (w_1183_, new_in6[2], w_1337_);
and (w_0026_, w_2051_, w_0829_);
nor (w_0369_, w_1644_, w_0830_);
nand (w_0877_, w_0985_, w_1140_);
and (w_0209_, w_1769_, w_0756_);
xor (w_1121_, w_1866_, w_0991_);
not (w_0932_, new_in6[2]);
and (w_1056_, new_in4[2], new_in1[0]);
nand (w_1179_, w_0726_, w_0583_);
xor (w_0807_, w_0752_, w_0630_);
nand (w_1787_, w_1322_, w_0303_);
nand (w_1945_, w_0511_, w_0125_);
xor (w_0746_, w_0218_, w_0059_);
xor (w_0217_, w_1071_, w_0144_);
or (w_1354_, w_1708_, w_1924_);
nand (w_1238_, w_1269_, w_1173_);
and (w_1471_, w_1147_, w_1614_);
not (w_0529_, new_in9[2]);
xor (w_0481_, w_0050_, w_1020_);
and (w_1973_, w_0085_, w_1745_);
nand (w_1374_, w_1548_, w_0297_);
and (w_0361_, w_1873_, w_1962_);
nand (w_1508_, w_0082_, w_0355_);
nand (w_1754_, w_1100_, w_0554_);
xor (w_1560_, new_in1[2], new_in3[5]);
nand (w_0335_, w_0372_, w_1011_);
nand (w_1779_, w_1380_, w_0877_);
nor (w_0804_, new_in10[1], new_in3[1]);
xor (w_1337_, new_in2[4], new_in5[5]);
nand (w_0437_, w_0347_, w_0573_);
nand (w_1632_, w_1946_, w_1817_);
nand (w_1069_, w_1318_, w_1268_);
xor (w_0870_, w_1519_, w_0337_);
xor (w_0112_, new_in6[4], w_0123_);
nand (w_1856_, w_0395_, w_0477_);
xor (w_0926_, w_1010_, w_1001_);
xor (w_1369_, w_1947_, w_0872_);
and (w_1649_, w_1857_, w_1563_);
xor (w_1415_, new_in8[3], w_0459_);
nand (w_1492_, w_1275_, w_1863_);
and (w_0230_, w_0177_, w_1387_);
xor (w_1036_, w_1038_, w_1468_);
and (w_1211_, new_in9[1], new_in1[1]);
and (w_0839_, w_0957_, w_2004_);
and (w_1405_, new_in8[4], new_in1[2]);
nand (w_1805_, w_0109_, w_1751_);
nand (w_1712_, w_0726_, w_1047_);
nand (w_1196_, w_0676_, w_1048_);
or (w_0600_, w_1707_, w_0420_);
and (w_1900_, new_in5[0], new_in8[0]);
xor (w_1168_, w_1613_, w_0457_);
nand (w_0704_, w_2071_, w_0389_);
and (w_1855_, w_2095_, w_1018_);
nand (w_0789_, w_1794_, w_0402_);
nand (w_0541_, w_1623_, w_0215_);
and (w_1647_, new_in10[0], new_in6[0]);
xor (w_0139_, new_in4[7], new_in6[3]);
nand (w_1247_, w_0726_, w_0401_);
nand (w_1227_, w_0088_, w_1775_);
xor (w_1684_, w_1861_, w_0146_);
xor (w_1355_, w_0952_, w_1569_);
or (w_0251_, w_0726_, w_1241_);
and (w_0601_, new_in8[3], new_in9[4]);
xor (w_1306_, w_0503_, w_1328_);
not (w_1426_, new_in6[0]);
or (w_1513_, w_1343_, w_0323_);
or (w_1275_, w_1693_, new_in6[7]);
xor (w_1063_, w_1517_, w_1272_);
xor (w_1236_, w_1725_, w_1891_);
xor (w_0816_, w_1302_, w_1245_);
or (w_1058_, w_0217_, w_2032_);
xor (w_0852_, w_0836_, w_0995_);
or (w_0152_, w_0200_, w_1122_);
or (w_1009_, w_1411_, w_1463_);
nand (w_0985_, w_0726_, w_0917_);
and (w_1326_, new_in2[6], new_in5[4]);
and (w_0578_, new_in9[6], new_in8[0]);
nand (w_0576_, w_1613_, w_0457_);
xor (w_1413_, w_0751_, w_0540_);
xor (w_0891_, w_0277_, w_1167_);
or (w_0957_, w_1755_, w_1082_);
xor (w_1731_, w_0250_, w_1540_);
xor (w_0233_, new_in6[3], w_0002_);
or (w_1184_, w_0726_, w_1504_);
or (w_1962_, w_0277_, w_1167_);
nand (w_0771_, new_in1[0], new_in8[6]);
xor (w_0297_, new_in11[0], w_1495_);
and (w_0946_, new_in8[0], new_in3[0]);
or (w_0163_, w_1708_, w_1171_);
xor (w_0184_, new_in6[7], w_0815_);
xor (w_0172_, w_0354_, w_1126_);
xor (w_0669_, new_in6[1], new_in11[0]);
and (w_1319_, w_0391_, w_0971_);
nand (w_1941_, w_1753_, w_1570_);
not (w_0040_, new_in2[4]);
xor (w_0424_, w_0741_, w_1113_);
xor (w_1927_, w_1523_, w_0955_);
nand (w_0765_, w_1857_, w_0546_);
nand (w_1668_, w_0019_, w_1445_);
nand (w_0474_, w_1237_, w_0415_);
nand (w_0592_, w_1708_, w_0883_);
nand (w_0005_, new_in1[0], new_in1[1]);
nand (w_0085_, w_1161_, new_in9[3]);
nand (w_0334_, w_1572_, w_1625_);
nand (w_0153_, w_1198_, w_1512_);
xor (w_1372_, new_in9[2], new_in1[1]);
nand (w_0377_, w_0319_, w_1945_);
xor (w_0519_, new_in3[1], w_2000_);
nand (w_1688_, w_0372_, w_1922_);
nand (w_0648_, w_1857_, w_1687_);
xor (w_1884_, new_in10[1], new_in3[2]);
xor (w_0907_, new_in10[3], new_in6[7]);
nand (w_1877_, new_in4[8], new_in8[6]);
and (w_1283_, new_in5[0], new_in2[3]);
nand (w_1494_, w_0200_, w_1604_);
and (w_1285_, new_in9[0], new_in8[0]);
xor (w_1686_, new_in9[3], new_in1[2]);
and (w_0210_, new_in9[2], new_in1[2]);
xor (w_1051_, new_in6[0], new_in8[6]);
xor (w_2061_, w_1949_, w_1288_);
nand (w_0225_, w_1708_, w_1461_);
nand (w_1987_, w_1857_, w_1709_);
not (w_1803_, new_in4[1]);
and (w_0486_, w_0939_, w_1537_);
nand (new_out9[3], w_0860_, w_0441_);
nand (w_1643_, w_1949_, w_1288_);
nand (w_1575_, w_0726_, w_1119_);
xor (w_0898_, w_1988_, w_1323_);
nand (w_2048_, w_0784_, w_0977_);
nand (w_1641_, w_0752_, w_0630_);
and (w_0378_, new_in8[3], new_in9[1]);
nand (w_1475_, w_1162_, w_0192_);
and (w_0952_, new_in5[1], new_in6[5]);
xor (w_1141_, w_1536_, w_0141_);
xor (w_1749_, new_in10[1], new_in4[1]);
xor (w_0410_, new_in5[3], w_0079_);
nand (w_2018_, w_1708_, w_0246_);
xor (w_0393_, new_in5[0], new_in2[1]);
nand (w_1173_, w_0787_, w_0831_);
xor (w_1408_, w_0482_, w_0825_);
and (w_0021_, new_in8[2], new_in11[0]);
or (w_1493_, w_0404_, w_2063_);
nand (w_1980_, w_0284_, w_0412_);
or (w_0214_, w_0200_, w_2014_);
and (w_1499_, new_in9[1], new_in8[5]);
nand (w_0886_, w_1708_, w_0264_);
nand (w_0375_, w_0331_, w_1231_);
xor (w_1589_, w_2093_, w_0881_);
xor (w_1148_, new_in9[4], new_in1[2]);
nand (w_1324_, new_in5[1], new_in2[1]);
xor (w_0150_, new_in5[2], w_0806_);
nand (w_1909_, w_1857_, w_1236_);
xor (w_0247_, w_0286_, w_1444_);
xor (w_1265_, w_0899_, w_0740_);
nand (w_0672_, w_0372_, w_0234_);
xor (w_1833_, new_in4[2], new_in6[2]);
nand (w_0485_, w_1291_, w_2092_);
xor (w_0188_, new_in11[1], w_0338_);
xor (w_0607_, w_0040_, new_in3[3]);
and (w_2001_, w_2010_, w_1714_);
xor (w_0916_, new_in3[1], w_0249_);
nand (w_1850_, w_1545_, new_in7[0]);
xor (w_1266_, w_0021_, w_1006_);
nand (w_0605_, w_0243_, w_0046_);
nand (w_1940_, w_1926_, w_0645_);
nand (w_1790_, w_0436_, w_1516_);
xor (w_0467_, w_1097_, w_1339_);
xor (w_1710_, w_0269_, w_0811_);
xor (w_1393_, w_2054_, w_1991_);
and (w_1610_, w_0826_, w_0912_);
and (w_1457_, w_2047_, w_1267_);
xor (w_0338_, new_in9[3], new_in9[4]);
nand (w_1143_, w_0217_, w_0743_);
nand (w_0403_, w_0932_, w_0862_);
nand (w_0215_, w_0609_, w_0111_);
nand (w_0413_, w_1536_, w_0141_);
and (w_1174_, new_in10[3], new_in6[2]);
nand (w_0259_, w_1708_, w_1446_);
xor (w_1988_, w_1283_, w_0292_);
and (w_0419_, new_in5[0], new_in1[0]);
and (w_1756_, w_1484_, w_0498_);
nand (w_0092_, w_1548_, w_1506_);
nand (w_1484_, new_in2[7], w_0193_);
xor (w_2081_, new_in1[2], new_in3[2]);
and (w_0950_, w_1677_, w_0627_);
or (w_0466_, w_0726_, w_1634_);
and (w_0252_, new_in8[2], new_in9[4]);
xor (w_0772_, w_0784_, w_0977_);
and (w_0882_, w_0556_, w_0444_);
and (w_2067_, w_1979_, w_1279_);
xor (w_0457_, new_in4[1], new_in8[1]);
nand (w_1485_, new_in11[0], new_in7[1]);
and (w_1054_, w_0741_, w_1373_);
xor (w_1164_, w_1921_, w_1145_);
nand (w_0525_, w_1133_, w_1037_);
xor (w_0244_, w_1042_, w_1165_);
nand (w_0274_, w_1081_, w_0961_);
nand (w_0499_, w_0970_, w_0616_);
and (w_1392_, w_0037_, w_1194_);
xor (w_1762_, w_0852_, w_2024_);
not (w_0492_, w_1648_);
not (w_0560_, new_in8[4]);
nand (w_1075_, w_0935_, w_1721_);
xor (w_1897_, w_1209_, w_0469_);
xor (w_0630_, new_in5[3], new_in2[3]);
and (w_0693_, w_0163_, w_0232_);
and (w_1071_, new_in11[0], new_in7[1]);
xor (w_1671_, new_in6[8], new_in2[3]);
nand (w_0318_, w_1857_, w_0999_);
xor (w_0032_, new_in2[7], new_in5[8]);
and (new_out8[0], w_0262_, w_0152_);
xor (w_0843_, w_1698_, w_0278_);
nand (w_2031_, w_0090_, w_2037_);
nand (w_2035_, w_0053_, w_0587_);
nand (w_0236_, w_1406_, new_in1[2]);
and (new_out5[0], w_1251_, w_0027_);
nand (w_0756_, w_1795_, w_0512_);
xor (w_0453_, w_1289_, w_1629_);
not (w_1252_, new_in8[2]);
xor (w_0566_, w_1012_, w_0055_);
xor (w_0940_, new_in2[7], w_0763_);
xor (w_0477_, w_0361_, w_0681_);
or (w_0640_, w_1967_, w_1931_);
nand (w_1483_, w_0305_, w_0374_);
nand (w_1367_, w_0200_, w_2062_);
nand (w_1573_, w_0726_, w_0738_);
nand (w_0532_, w_0726_, w_1234_);
and (w_0006_, w_1426_, new_in4[0]);
nand (w_0927_, w_1708_, w_1787_);
not (w_0755_, new_in2[7]);
xor (w_1682_, new_in9[5], new_in1[3]);
nand (w_1866_, w_1477_, w_1314_);
xor (w_1574_, w_0637_, w_1372_);
or (w_0290_, w_0726_, w_0705_);
and (w_0089_, w_0217_, w_1772_);
nand (w_1862_, w_0637_, w_1372_);
and (w_0020_, w_0217_, w_1712_);
not (w_0505_, new_in4[4]);
or (w_1559_, new_in10[0], new_in3[0]);
nand (w_0402_, w_1976_, w_1336_);
xor (w_0938_, w_0271_, w_0426_);
and (w_0976_, new_in9[2], w_0162_);
or (w_1658_, w_1381_, w_1995_);
nand (w_0587_, w_0217_, w_0213_);
nand (w_0169_, w_0979_, w_0589_);
nand (w_1436_, w_0354_, w_1126_);
and (w_1672_, w_0069_, w_1996_);
xor (w_0064_, w_1586_, w_1558_);
xor (w_0117_, new_in6[3], w_0506_);
xor (w_0706_, new_in5[0], new_in5[1]);
nand (w_1794_, new_in10[3], new_in4[3]);
or (w_0306_, w_0200_, w_0462_);
or (w_0959_, w_0904_, w_0793_);
xor (w_1347_, new_in9[0], new_in1[3]);
nand (w_1032_, w_1781_, w_0004_);
xor (w_0925_, w_0962_, w_1998_);
not (w_1042_, new_in4[2]);
xor (w_0367_, w_0384_, w_0304_);
xor (w_1934_, new_in10[3], w_1528_);
or (w_1930_, w_0962_, w_0369_);
xor (w_0812_, w_1001_, w_0420_);
nand (w_1977_, w_0174_, w_1819_);
nand (w_1078_, w_1072_, w_0198_);
xor (w_1014_, w_1356_, w_0095_);
nand (w_0892_, w_0217_, w_1980_);
and (w_2095_, new_in1[0], new_in3[0]);
and (w_0609_, new_in3[0], w_1129_);
xor (w_1539_, w_0035_, w_1762_);
and (w_1470_, w_1764_, w_1311_);
and (w_0698_, w_0726_, w_1044_);
and (w_0563_, w_1639_, w_0841_);
xor (w_1598_, new_in6[0], w_1999_);
xor (w_0226_, new_in2[2], new_in5[3]);
xor (w_1898_, new_in10[1], new_in4[0]);
xor (w_0100_, w_1025_, w_0624_);
or (w_1750_, w_0301_, w_0221_);
xor (w_1323_, w_0116_, w_0661_);
nand (w_0347_, w_0782_, w_1720_);
or (w_0231_, w_0217_, w_1502_);
nor (w_1995_, w_0114_, new_in1[0]);
xor (w_0307_, new_in1[3], w_1818_);
nand (w_0025_, w_1337_, w_0289_);
xor (w_1872_, new_in6[5], new_in7[0]);
xor (w_1018_, new_in1[1], new_in3[1]);
nand (w_0250_, w_1864_, w_0966_);
xor (w_0622_, w_0030_, w_1703_);
and (w_0559_, w_1921_, new_in4[5]);
xor (w_1654_, w_1288_, w_0895_);
xor (w_0108_, w_1301_, w_0320_);
xor (w_0344_, w_0381_, w_0072_);
xor (w_0817_, w_0630_, w_2058_);
and (w_1417_, new_in8[2], w_0291_);
xor (w_1557_, w_1967_, new_in8[0]);
nand (w_1679_, w_1478_, w_1149_);
xor (w_0312_, w_0714_, w_0770_);
xor (w_0846_, new_in11[1], new_in7[1]);
xor (w_0853_, w_0787_, w_0831_);
and (w_0142_, new_in9[3], new_in9[4]);
nand (w_1860_, w_0501_, w_0778_);
xor (w_0633_, new_in8[4], new_in9[4]);
xor (w_1984_, new_in4[6], new_in6[2]);
nand (w_1335_, w_0168_, w_0851_);
xor (w_1619_, w_0725_, w_1120_);
xor (w_0267_, new_in3[2], w_1682_);
xor (w_1430_, w_1814_, w_1378_);
nand (w_2052_, w_0726_, w_1164_);
and (w_1435_, w_0121_, w_0538_);
and (w_1128_, new_in10[3], new_in7[0]);
nand (w_1085_, w_1521_, w_1442_);
xor (w_1122_, w_2010_, w_1714_);
xor (w_1700_, w_1587_, w_0103_);
xor (w_0038_, w_1431_, w_1160_);
nand (w_0204_, w_0790_, w_1662_);
xor (w_1234_, w_2011_, w_1238_);
or (w_0158_, w_1192_, w_1451_);
nand (w_1907_, new_in11[1], w_0783_);
xor (w_0122_, w_1357_, w_0219_);
nand (w_1646_, w_0121_, w_0538_);
xor (w_0543_, w_0827_, new_in4[3]);
xor (w_1451_, new_in9[1], w_0260_);
nand (new_out6[1], w_1135_, w_0275_);
nand (w_0364_, w_1429_, w_1741_);
xor (w_2026_, w_2064_, w_0155_);
xor (w_1563_, w_1985_, w_1655_);
xor (w_0508_, w_0395_, w_1656_);
nand (w_0978_, new_in2[4], new_in5[5]);
nor (w_0298_, w_0408_, w_0289_);
xor (w_1116_, w_0770_, w_1224_);
nand (w_1895_, w_0335_, w_2098_);
nand (w_1838_, w_1857_, w_1735_);
and (w_0353_, w_0022_, w_0413_);
xor (w_1139_, w_1157_, w_1095_);
nand (w_0133_, w_1921_, w_1337_);
xor (w_0889_, new_in3[6], w_1791_);
xor (w_0183_, w_1521_, w_1442_);
xor (w_0581_, w_1892_, w_0117_);
xor (w_0161_, w_1115_, w_0748_);
or (w_1990_, w_0217_, w_1601_);
xor (w_1241_, w_0847_, w_0209_);
nand (w_1084_, w_1548_, w_0692_);
and (w_1156_, new_in10[3], new_in2[1]);
xor (w_1246_, w_1104_, w_1466_);
xor (w_1255_, new_in6[2], w_0862_);
xor (w_0261_, w_0862_, w_0514_);
xor (w_0110_, w_1519_, w_1582_);
nand (w_0670_, w_1548_, w_0281_);
nand (w_0387_, w_0265_, w_1178_);
or (w_1099_, w_0726_, w_1448_);
nand (w_0270_, new_in2[0], w_0852_);
xor (w_1801_, w_1187_, w_0113_);
and (w_0980_, new_in10[2], new_in2[0]);
nand (w_0280_, w_1718_, w_0574_);
nand (w_0820_, w_0919_, w_0307_);
nand (w_0972_, w_0857_, w_0236_);
nand (new_out1[3], w_1757_, w_1809_);
and (w_1416_, w_0287_, w_0071_);
or (w_0649_, w_1031_, w_1489_);
nand (w_1123_, w_1509_, w_0593_);
xor (w_1172_, w_1217_, w_0188_);
xor (w_0757_, w_0621_, w_1500_);
nor (w_0086_, w_0784_, w_0674_);
xor (w_1882_, w_0889_, w_1675_);
nand (w_1915_, w_0843_, w_0261_);
or (w_1617_, w_0361_, w_0681_);
nor (w_0987_, new_in6[0], new_in4[0]);
xor (w_0000_, w_1668_, w_0351_);
xor (w_1385_, w_0511_, w_0125_);
xor (w_1026_, w_0686_, w_1870_);
and (w_1082_, w_1658_, w_0803_);
nand (new_out10[3], w_0434_, w_1954_);
xor (w_1092_, w_1252_, w_0852_);
and (w_1212_, w_0741_, w_0753_);
nand (w_0345_, w_1366_, w_1968_);
xor (w_1465_, w_0046_, w_0244_);
nand (w_0484_, w_0513_, new_in5[6]);
and (w_0725_, w_0973_, w_0762_);
xor (w_1250_, w_0252_, w_0518_);
xor (w_0844_, w_2081_, w_1168_);
and (w_1159_, w_0385_, w_2031_);
or (w_1906_, w_0200_, w_0034_);
xor (w_1664_, w_0654_, w_0440_);
nand (w_1294_, w_0510_, w_1871_);
nand (w_1472_, w_0453_, w_1957_);
xor (w_0301_, w_0565_, w_2006_);
nand (w_0691_, w_2078_, w_0646_);
not (w_1406_, new_in1[1]);
nand (w_0526_, w_0217_, w_0744_);
nand (w_1780_, w_0520_, w_0178_);
nor (w_0703_, new_in9[1], new_in8[1]);
xor (w_2023_, new_in10[0], new_in3[3]);
nand (w_0567_, w_0708_, w_0855_);
xor (w_1763_, w_1882_, w_0324_);
or (w_1158_, w_0503_, w_1328_);
xor (w_0697_, w_0485_, w_1501_);
nand (w_1008_, w_1630_, new_in9[2]);
xor (w_1244_, new_in10[2], new_in4[2]);
nand (w_1304_, w_0175_, w_1621_);
nand (w_0264_, w_0590_, w_1786_);
xor (w_0865_, w_1776_, w_0456_);
xor (w_1476_, w_0070_, w_1347_);
or (w_1190_, w_1708_, w_1607_);
nand (w_0822_, w_1252_, new_in9[1]);
xor (w_1946_, w_1839_, w_0407_);
xor (w_2024_, w_1060_, w_1130_);
xor (w_1163_, w_0007_, w_0754_);
xor (w_1053_, w_0419_, w_1474_);
not (w_1338_, w_1519_);
nand (w_0826_, new_in9[2], w_0273_);
and (w_0324_, w_0044_, w_1737_);
nand (w_0208_, w_0217_, w_1851_);
nand (w_1944_, w_0217_, w_1692_);
nand (new_out6[3], w_1807_, w_0653_);
not (w_1967_, new_in5[0]);
xor (w_1924_, w_1760_, w_1690_);
nand (w_2057_, w_1708_, w_1868_);
not (w_1287_, w_1288_);
not (w_0878_, new_in9[4]);
and (w_1810_, new_in6[0], new_in4[0]);
xor (w_0321_, w_0046_, w_0807_);
or (w_0322_, w_0123_, w_1577_);
xor (w_0955_, w_1936_, w_1820_);
not (w_1025_, w_1681_);
and (w_1514_, w_1853_, w_0814_);
xor (w_0125_, new_in3[1], new_in2[2]);
xor (w_0700_, w_0921_, w_1180_);
and (w_0751_, new_in9[0], new_in1[3]);
or (w_0181_, w_1883_, w_1686_);
xor (w_0281_, w_0964_, w_1185_);
nand (w_2074_, w_0375_, w_1987_);
not (w_1548_, w_0726_);
or (w_0558_, w_1684_, w_0452_);
xor (w_1463_, w_1288_, w_2038_);
xor (w_2007_, w_1348_, w_0948_);
and (w_1795_, new_in11[0], w_1495_);
xor (w_0194_, w_0145_, w_2066_);
nand (w_1812_, new_in1[3], w_1818_);
or (w_0690_, w_0755_, new_in6[3]);
nand (w_2013_, w_0067_, new_in5[7]);
or (w_0824_, w_0200_, w_0400_);
xor (w_1953_, new_in4[6], w_0674_);
nand (w_1419_, w_0726_, w_2091_);
nand (w_1543_, w_1573_, w_0875_);
nand (w_0037_, new_in6[7], new_in2[2]);
xor (w_0715_, new_in10[2], w_0582_);
not (w_1434_, w_1357_);
xor (w_1799_, new_in1[0], w_0818_);
and (w_1195_, new_in10[3], new_in2[0]);
nand (w_0900_, w_1834_, w_1773_);
or (w_1551_, w_1930_, w_0571_);
or (w_0254_, w_0248_, w_1628_);
nand (w_1207_, w_1708_, w_1824_);
xor (w_1870_, w_1392_, w_1671_);
and (w_1034_, w_0600_, w_0934_);
nand (w_0228_, w_0168_, w_1036_);
xor (w_0383_, w_0075_, w_0074_);
xor (w_0171_, new_in3[2], w_1093_);
or (w_1409_, w_0559_, w_1984_);
xor (w_0665_, w_1261_, w_0543_);
xor (w_2092_, new_in10[3], new_in7[0]);
xor (w_2010_, new_in10[0], new_in9[2]);
nand (w_1802_, new_in10[3], new_in4[2]);
and (w_1013_, w_2088_, w_0008_);
xor (w_2082_, w_0628_, w_1172_);
nand (w_2022_, new_in1[2], new_in3[3]);
nand (w_1785_, new_in3[2], new_in2[2]);
nand (w_1845_, w_1800_, w_0905_);
nand (w_1696_, w_0864_, w_1346_);
xor (w_0068_, w_1146_, w_0491_);
xor (w_1232_, w_1016_, w_1733_);
and (w_0702_, new_in10[1], new_in2[0]);
nand (w_0589_, w_0021_, w_1006_);
nand (w_0099_, new_in4[1], new_in8[1]);
xor (w_0683_, w_0505_, new_in10[5]);
nand (w_1865_, w_0168_, w_1898_);
or (w_1532_, w_0726_, w_0253_);
nand (w_1223_, w_0168_, w_0712_);
and (w_0429_, new_in1[1], new_in8[5]);
xor (w_1561_, w_0449_, w_0950_);
xor (w_0066_, w_1406_, w_1598_);
nand (w_0399_, w_1324_, w_0093_);
nor (w_1965_, w_1789_, w_1327_);
and (w_1166_, new_in4[0], w_1326_);
xor (w_1587_, w_0567_, w_0781_);
xor (w_0675_, new_in8[1], new_in11[1]);
nand (w_0348_, w_1857_, w_0370_);
nand (w_1221_, w_1318_, w_1218_);
nand (w_0887_, w_0726_, w_0853_);
nand (w_2019_, w_0882_, w_1407_);
nand (w_1771_, w_1673_, w_1404_);
nand (w_1723_, w_0636_, w_0387_);
and (w_1425_, w_1857_, w_1524_);
nand (w_0667_, w_0765_, w_1680_);
nand (w_1948_, w_1857_, w_1265_);
xor (w_0072_, new_in4[2], new_in1[0]);
nand (w_0294_, w_0862_, w_0101_);
and (w_1625_, w_1915_, w_0212_);
nand (w_1424_, w_1857_, w_1121_);
nand (w_0391_, w_0852_, w_2024_);
xor (w_0689_, new_in8[2], new_in9[1]);
xor (w_0380_, w_1068_, w_0226_);
nand (w_0873_, new_in5[8], new_in3[5]);
and (w_0023_, w_0861_, w_0679_);
nand (w_1919_, w_0257_, w_2057_);
nand (w_1481_, w_0217_, w_1487_);
nand (w_0392_, w_0217_, w_1566_);
and (w_0135_, w_1708_, w_1197_);
nand (w_1489_, w_0439_, w_1907_);
nand (w_0268_, w_0377_, w_0042_);
nand (new_out9[0], w_1274_, w_0300_);
nand (w_1969_, w_0488_, new_in6[6]);
nand (w_1645_, w_1209_, w_0469_);
nand (w_0327_, w_1729_, w_0772_);
nand (w_0996_, w_1648_, w_1222_);
nand (w_1165_, w_0350_, w_1899_);
xor (w_1804_, w_1021_, w_2011_);
nor (w_1923_, w_0040_, new_in5[5]);
xor (w_0050_, w_1112_, w_0126_);
and (w_1843_, w_0217_, w_1836_);
and (new_out8[2], w_0147_, w_0306_);
and (w_0007_, new_in6[5], new_in7[0]);
nand (w_1363_, w_1776_, w_0456_);
nand (new_out7[1], w_0084_, w_0673_);
or (w_1972_, w_0200_, w_0643_);
xor (w_0620_, new_in10[3], new_in9[3]);
nand (w_1482_, w_1862_, w_0866_);
nand (w_0854_, w_1023_, w_0259_);
and (w_1768_, w_1428_, w_1341_);
xor (w_1638_, w_0317_, w_1695_);
xor (w_1721_, w_1546_, w_0909_);
or (w_1853_, w_1708_, w_1626_);
xor (w_0920_, new_in1[0], w_1385_);
and (w_0523_, w_2048_, w_0327_);
xor (w_1124_, w_1029_, w_0227_);
xor (w_0134_, new_in4[0], new_in2[4]);
nand (w_1896_, new_in4[7], new_in8[5]);
nand (w_0829_, w_0725_, w_1120_);
and (w_1328_, w_0390_, w_0822_);
and (w_1594_, w_0180_, w_0602_);
nor (w_0144_, new_in9[2], new_in1[3]);
xor (w_0833_, w_0689_, w_1741_);
xor (w_0001_, w_1999_, w_0732_);
nand (w_0879_, w_0774_, w_0516_);
nand (w_1537_, w_1708_, w_0105_);
or (w_0874_, w_0726_, w_1700_);
nand (w_1382_, w_1708_, w_1790_);
or (w_0396_, w_0200_, w_0508_);
xor (w_1874_, w_0017_, w_2080_);
nand (w_1040_, w_1548_, w_0417_);
xor (w_1653_, new_in6[3], w_0123_);
xor (w_1224_, w_1879_, w_1810_);
and (w_1033_, w_1289_, w_1629_);
nand (w_0552_, new_in1[3], new_in3[3]);
and (w_2080_, w_0332_, w_1507_);
nand (w_0777_, w_1828_, w_2077_);
nor (w_0888_, w_0082_, w_0703_);
and (w_0522_, w_0239_, w_0980_);
xor (w_0473_, w_1435_, w_1114_);
xor (w_1048_, new_in10[2], new_in3[5]);
not (w_1021_, w_0258_);
and (w_1193_, w_1545_, w_2022_);
nand (w_0911_, w_0217_, w_0065_);
xor (w_1079_, w_2028_, w_0238_);
nand (w_2004_, w_0529_, new_in1[2]);
nand (w_1240_, w_0129_, w_1191_);
nand (w_1387_, w_1151_, w_1465_);
xor (w_1528_, w_1594_, w_0112_);
or (w_0553_, w_1110_, w_1260_);
and (w_0340_, w_1286_, w_1830_);
nand (w_1377_, new_in8[4], w_0169_);
and (w_1478_, w_0128_, w_1049_);
nand (w_1086_, w_0023_, w_1250_);
and (w_2039_, w_1001_, w_0393_);
xor (w_1101_, w_1291_, w_2092_);
and (w_1330_, w_1708_, w_0231_);
nand (w_0517_, new_in10[1], w_1542_);
nand (w_0343_, w_1857_, w_1202_);
nand (w_0265_, w_1128_, w_0494_);
xor (w_0330_, w_1086_, w_1711_);
xor (w_0400_, new_in5[0], w_0987_);
nand (w_1073_, w_0662_, w_0597_);
nand (new_out4, w_1742_, w_0091_);
nand (w_1960_, new_in6[7], w_0815_);
nand (w_0677_, w_0200_, w_1580_);
or (w_0682_, w_0487_, w_1255_);
nand (w_0564_, w_0726_, w_0061_);
nand (w_1844_, w_1708_, w_1206_);
xor (w_1125_, new_in10[1], w_1139_);
and (w_1618_, w_0421_, w_0535_);
xor (w_1394_, new_in1[2], w_1063_);
xor (w_0061_, w_1151_, w_1465_);
nand (w_0863_, w_0372_, w_0611_);
nand (w_0979_, new_in8[3], new_in11[1]);
nand (w_1427_, w_0726_, w_1046_);
nand (w_1379_, new_in8[2], w_0852_);
or (w_0934_, w_0899_, w_0740_);
nand (w_0246_, w_1579_, w_0998_);
not (w_0770_, w_1001_);
nand (w_1816_, w_0871_, w_0268_);
xor (w_0730_, w_0837_, w_0579_);
xor (w_1352_, new_in4[3], new_in1[1]);
nand (w_1396_, w_0726_, w_1125_);
nand (w_1718_, w_0372_, w_1004_);
nand (w_0717_, new_in9[1], new_in1[4]);
and (w_0763_, w_0097_, w_1032_);
xor (w_0401_, w_1192_, w_1451_);
nand (w_1873_, w_1161_, new_in9[1]);
and (w_0964_, w_0316_, w_0254_);
xor (w_0317_, w_0984_, w_0689_);
nand (w_1115_, w_1201_, w_0012_);
or (w_1681_, w_0325_, w_0963_);
xor (w_0862_, new_in2[5], new_in5[6]);
xor (w_0616_, new_in4[3], new_in10[4]);
nand (new_out9[2], w_1590_, w_1389_);
nand (w_0331_, w_0726_, w_1934_);
xor (w_0988_, new_in4[1], new_in3[2]);
xor (w_1253_, w_1636_, w_0652_);
nand (w_1729_, w_1508_, w_1771_);
xor (w_1145_, new_in10[0], w_1447_);
and (w_2044_, new_in10[5], w_1703_);
nand (w_1089_, new_in8[1], new_in7[1]);
or (w_1370_, w_1155_, w_1822_);
and (w_0613_, w_0381_, w_2060_);
nand (w_1488_, w_1338_, w_1582_);
nand (w_1360_, new_in10[4], new_in7[1]);
nand (w_0660_, w_0168_, w_0157_);
xor (w_1530_, w_1390_, w_1503_);
and (w_0963_, w_1300_, w_1905_);
nand (w_1536_, w_1739_, w_1854_);
xor (w_2037_, new_in8[1], w_1373_);
nand (w_1242_, w_0694_, w_0718_);
nand (w_1775_, w_1599_, w_0675_);
or (w_1072_, w_1708_, w_1850_);
nand (w_1611_, w_1230_, w_0057_);
nand (w_2016_, w_1879_, w_0006_);
nand (w_0394_, w_1857_, w_0812_);
xor (w_0584_, w_2028_, w_0907_);
xor (w_0503_, new_in8[3], new_in9[2]);
nand (w_1038_, w_0496_, w_1085_);
and (w_1441_, new_in1[0], new_in3[2]);
nand (w_0922_, w_0200_, w_0486_);
nand (w_0997_, w_0933_, w_1526_);
xor (w_0469_, w_1916_, w_1079_);
nand (w_0760_, w_1705_, w_2065_);
xor (w_1407_, w_0453_, w_1957_);
nand (w_0733_, w_2083_, w_0431_);
nand (w_0329_, w_0211_, w_0903_);
nand (w_1890_, new_in8[3], new_in4[5]);
or (w_1858_, w_0545_, w_0285_);
xor (w_0783_, new_in1[0], new_in3[1]);
and (w_1411_, w_0958_, w_0366_);
xor (w_1848_, w_1088_, w_0727_);
nand (w_1280_, new_in2[5], new_in5[3]);
nand (w_1609_, w_1879_, w_0737_);
xor (w_0685_, w_1174_, w_0314_);
nand (w_0617_, w_0726_, w_0256_);
nand (w_1395_, w_0160_, w_0610_);
or (w_1739_, w_1530_, w_2089_);
nand (w_1992_, w_1744_, w_1040_);
or (w_1517_, new_in10[3], new_in3[3]);
or (w_1226_, w_0964_, w_1185_);
xor (w_1512_, w_0210_, w_0000_);
xor (w_0507_, w_0938_, w_1383_);
nor (w_0323_, w_1373_, w_0399_);
xor (w_0405_, w_1666_, w_0340_);
and (w_0079_, w_0470_, w_0893_);
xor (w_0593_, w_0551_, w_0032_);
xor (w_0686_, w_0471_, w_1966_);
or (w_1867_, w_1425_, w_0835_);
and (w_0621_, w_0060_, w_0158_);
or (w_0379_, w_0862_, w_2021_);
xor (w_1975_, w_0393_, w_1045_);
xor (w_2027_, new_in11[0], new_in9[3]);
nand (w_1362_, new_in2[5], new_in5[1]);
xor (w_0572_, w_0381_, w_1258_);
xor (w_1468_, w_1050_, w_0537_);
xor (w_0918_, new_in4[7], w_2034_);
and (w_0360_, new_in6[5], new_in2[0]);
not (w_2060_, w_0072_);
nand (w_0197_, w_0819_, w_2079_);
nand (w_0735_, w_0308_, w_1541_);
and (w_1343_, w_1373_, w_0399_);
xor (w_1291_, w_1108_, w_1290_);
nand (w_1704_, w_1364_, w_1556_);
nand (w_2070_, w_1990_, w_1747_);
xor (w_0680_, new_in1[0], new_in1[1]);
xor (w_0748_, new_in4[2], new_in3[3]);
and (w_1296_, w_1916_, w_1079_);
xor (w_2077_, new_in10[3], new_in4[2]);
and (w_0062_, new_in10[2], w_1903_);
nand (w_0910_, w_1708_, w_1583_);
xor (w_1793_, w_0367_, w_0891_);
xor (w_0017_, w_1499_, w_0858_);
nand (w_0639_, w_0726_, w_1443_);
nand (new_out6[2], w_1606_, w_0228_);
xor (w_1031_, w_0689_, w_1917_);
xor (w_1982_, w_0248_, w_1628_);
and (w_0463_, new_in8[0], new_in7[0]);
nor (w_1496_, w_0217_, w_0321_);
xor (w_1554_, w_2066_, w_0669_);
and (w_1300_, new_in1[0], new_in3[1]);
nand (w_0262_, w_0200_, w_1768_);
xor (w_0981_, new_in9[5], new_in1[4]);
nand (w_1281_, w_0250_, w_1540_);
xor (w_1447_, w_0862_, w_1923_);
nand (w_1796_, new_in8[2], new_in9[1]);
xor (w_2072_, new_in11[0], w_0785_);
nand (w_0175_, w_1584_, w_1176_);
nand (w_1286_, new_in9[3], w_1293_);
nand (w_1199_, w_1075_, w_1005_);
and (new_out1[1], w_0423_, w_0214_);
or (w_1178_, w_1128_, w_0494_);
xor (w_0138_, w_0299_, w_1136_);
xor (w_1310_, new_in1[1], w_0773_);
xor (w_0766_, w_1927_, w_1224_);
xor (w_0901_, w_1781_, w_0004_);
or (w_1620_, w_0200_, w_1101_);
xor (w_1656_, w_0054_, w_0124_);
nand (w_0787_, w_1609_, w_1534_);
xor (w_0432_, w_0094_, w_0365_);
xor (w_1777_, w_1435_, w_0848_);
or (w_0728_, w_0726_, w_0272_);
xor (w_0806_, new_in1[3], new_in3[6]);
not (w_0827_, new_in8[3]);
xor (w_1399_, new_in9[5], new_in9[4]);
nand (w_0016_, w_0200_, w_0416_);
xor (w_0055_, new_in1[6], w_1204_);
or (w_1050_, new_in4[2], new_in6[2]);
nand (w_0098_, w_0726_, w_0233_);
nand (w_0913_, new_in6[4], w_0505_);
and (w_1308_, w_0217_, w_0974_);
or (w_0255_, w_1181_, w_0846_);
nand (w_0176_, w_0168_, w_0697_);
xor (w_0465_, w_2033_, w_1806_);
nand (w_0619_, w_0217_, w_1552_);
xor (w_1711_, w_1321_, w_1219_);
nand (w_0764_, w_0217_, w_1992_);
xor (w_1825_, new_in4[6], new_in6[6]);
nor (w_1497_, w_0631_, w_0086_);
nand (w_1914_, w_0372_, w_0572_);
and (new_out11[1], w_0200_, w_1902_);
xor (w_1065_, w_1477_, w_1314_);
xor (w_1454_, new_in8[5], w_1777_);
or (w_0151_, w_0217_, w_1574_);
or (w_1043_, w_1103_, w_0193_);
xor (w_0937_, w_0352_, new_in8[6]);
nand (w_1400_, w_0726_, w_0757_);
nand (w_0315_, w_1548_, w_0245_);
xor (w_0645_, w_1310_, w_1403_);
and (w_0289_, w_1823_, w_1999_);
xor (w_1600_, w_0817_, w_0918_);
or (w_1218_, new_in4[3], new_in5[7]);
nand (w_1350_, new_in8[3], new_in9[0]);
nand (w_0041_, w_0372_, w_1619_);
and (w_0949_, w_0792_, w_1971_);
xor (w_1697_, w_0123_, w_0311_);
and (w_1673_, w_1285_, w_1792_);
and (w_1776_, new_in11[0], w_0701_);
nand (w_0524_, w_0200_, w_0931_);
and (w_0652_, new_in9[5], new_in8[2]);
or (w_1937_, w_1708_, w_1080_);
xor (w_1317_, w_0827_, w_1618_);
not (w_0067_, new_in2[6]);
nand (w_1566_, w_0164_, w_0290_);
xor (w_2064_, w_0656_, w_0283_);
xor (w_1901_, w_1661_, w_1309_);
nand (new_out10[0], w_0677_, w_1620_);
xor (w_0351_, w_1375_, w_0139_);
nand (w_0939_, w_0372_, w_1035_);
nand (w_1571_, w_1887_, w_0473_);
nand (w_1531_, w_0168_, w_0519_);
xor (w_1670_, w_0558_, w_1801_);
xor (w_1288_, w_2095_, w_1018_);
xor (w_2049_, w_0559_, w_1984_);
or (w_1097_, new_in9[5], new_in1[2]);
or (w_0087_, w_0200_, w_1849_);
nand (w_0992_, w_0372_, w_0502_);
and (new_out11[0], w_0200_, w_0115_);
xor (w_1510_, new_in2[7], new_in6[3]);
not (w_0114_, new_in9[0]);
xor (w_1572_, w_1124_, w_1697_);
nand (w_0179_, w_0168_, w_1479_);
nand (w_0726_, w_1458_, w_1576_);
nand (w_1024_, w_1708_, w_1779_);
xor (w_0738_, w_1931_, w_1233_);
nand (w_0275_, w_0168_, w_0183_);
or (w_0535_, w_0295_, w_1457_);
nand (w_0774_, new_in2[5], w_1803_);
or (w_1458_, w_0940_, w_1216_);
nand (w_0740_, w_0600_, w_1549_);
nor (w_1444_, new_in6[1], new_in4[5]);
and (w_1366_, w_1001_, w_1559_);
nand (w_0332_, w_1000_, w_0928_);
nand (w_1823_, w_0293_, w_1722_);
or (w_0326_, new_in6[3], new_in4[3]);
xor (w_1080_, w_1252_, w_1300_);
nand (w_1318_, new_in4[3], new_in5[7]);
or (w_1764_, w_1050_, w_0537_);
xor (w_1726_, w_1530_, w_2089_);
nand (w_0539_, new_in10[1], new_in4[1]);
xor (w_0650_, w_0722_, w_1859_);
xor (w_1113_, new_in10[2], new_in6[6]);
nand (w_0200_, w_1123_, w_1270_);
xor (w_1957_, new_in6[6], new_in3[1]);
and (w_1652_, w_0325_, w_1728_);
xor (w_0124_, new_in5[1], w_1560_);
nand (w_0845_, w_0726_, w_1920_);
xor (w_0111_, new_in3[1], w_1148_);
nand (w_1256_, w_0372_, w_1638_);
nand (w_0856_, w_0116_, w_0661_);
and (w_0800_, w_1503_, w_0634_);
and (w_1651_, w_0364_, w_1880_);
xor (w_0557_, w_0127_, w_0753_);
xor (w_0119_, w_1435_, w_1581_);
xor (w_1187_, w_0839_, w_0834_);
nand (w_0493_, w_0447_, w_1986_);
nand (w_0821_, w_0380_, w_1804_);
xor (w_1169_, new_in1[2], new_in5[2]);
xor (w_1129_, new_in9[3], new_in1[1]);
xor (w_1098_, w_1262_, w_1319_);
nand (w_0363_, w_0960_, w_0448_);
nand (w_0671_, w_2054_, w_1991_);
nand (w_2043_, w_0334_, w_0698_);
nor (w_1964_, w_1727_, w_1701_);
and (w_0120_, new_in9[5], new_in8[1]);
nand (w_0501_, w_0123_, w_1073_);
xor (w_1607_, w_0383_, w_0222_);
or (w_0890_, w_1708_, w_2072_);
xor (w_1727_, new_in5[2], new_in2[3]);
and (w_0598_, w_0378_, w_0550_);
nand (w_0883_, w_1522_, w_1538_);
endmodule
