module top_module (
    input wire  [2:0] in1_sub_module1,
    input wire  [2:0] in2_sub_module1,
    input wire  [2:0] in3_sub_module1,
    output wire [2:0] out1_sub_module1,
    output wire [2:0] out2_sub_module1,
    input wire  [2:0] in1_sub_module2,
    input wire  [2:0] in2_sub_module2,
    input wire  [2:0] in3_sub_module2,
    input wire  [2:0] in4_sub_module2,
    input wire  [2:0] in5_sub_module2,
    input wire  [2:0] in6_sub_module2,
    input wire  [2:0] in7_sub_module2,
    input wire  [2:0] in8_sub_module2,
    input wire  [2:0] in9_sub_module2,
    input wire  [2:0] in10_sub_module2,
    input wire  [2:0] in11_sub_module2,
    input wire  [2:0] in12_sub_module2,
    output wire [2:0] out1_sub_module2,
    output wire [2:0] out2_sub_module2,
    output wire [2:0] out3_sub_module2,
    output wire [2:0] out4_sub_module2,
    output wire [2:0] out5_sub_module2,
    output wire [2:0] out6_sub_module2,
    input wire  [8:0] in1_sub_module3,
    input wire  [8:0] in2_sub_module3,
    input wire  [8:0] in3_sub_module3,
    input wire  [8:0] in4_sub_module3,
    input wire  [6:0] in5_sub_module3,
    input wire  [6:0] in6_sub_module3,
    input wire  [6:0] in7_sub_module3,
    input wire  [6:0] in8_sub_module3,
    input wire  [6:0] in9_sub_module3,
    input wire  [1:0] in10_sub_module3,
    input wire  [1:0] in11_sub_module3,
    output wire       out1_sub_module3,
    output wire       out2_sub_module3,
    output wire [3:0] out3_sub_module3,
    output wire [3:0] out4_sub_module3,
    output wire [3:0] out5_sub_module3,
    output wire [3:0] out6_sub_module3,
    output wire [3:0] out7_sub_module3,
    output wire [3:0] out8_sub_module3,
    output wire [3:0] out9_sub_module3,
    output wire [3:0] out10_sub_module3,
    output wire [3:0] out11_sub_module3
);
    sub_module1 U1 (
        .in1(in1_sub_module1),
        .in2(in2_sub_module1),
        .in3(in3_sub_module1),
        .out1(out1_sub_module1),
        .out2(out2_sub_module1)
    );

    sub_module2 U2 (
        .in1(in1_sub_module2),
        .in2(in2_sub_module2),
        .in3(in3_sub_module2),
        .in4(in4_sub_module2),
        .in5(in5_sub_module2),
        .in6(in6_sub_module2),
        .in7(in7_sub_module2),
        .in8(in8_sub_module2),
        .in9(in9_sub_module2),
        .in10(in10_sub_module2),
        .in11(in11_sub_module2),
        .in12(in12_sub_module2),
        .out1(out1_sub_module2),
        .out2(out2_sub_module2),
        .out3(out3_sub_module2),
        .out4(out4_sub_module2),
        .out5(out5_sub_module2),
        .out6(out6_sub_module2)
    );

    sub_module3 U3 (
        .in1(in1_sub_module3),
        .in2(in2_sub_module3),
        .in3(in3_sub_module3),
        .in4(in4_sub_module3),
        .in5(in5_sub_module3),
        .in6(in6_sub_module3),
        .in7(in7_sub_module3),
        .in8(in8_sub_module3),
        .in9(in9_sub_module3),
        .in10(in10_sub_module3),
        .in11(in11_sub_module3),
        .out1(out1_sub_module3),
        .out2(out2_sub_module3),
        .out3(out3_sub_module3),
        .out4(out4_sub_module3),
        .out5(out5_sub_module3),
        .out6(out6_sub_module3),
        .out7(out7_sub_module3),
        .out8(out8_sub_module3),
        .out9(out9_sub_module3),
        .out10(out10_sub_module3),
        .out11(out11_sub_module3)
    );

endmodule
